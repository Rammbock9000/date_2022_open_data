--------------------------------------------------------------------------------
--                         ModuloCounter_64_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity ModuloCounter_64_component is
   port ( clk, rst : in std_logic;
          Counter_out : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of ModuloCounter_64_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk,rst)
	 variable count : std_logic_vector(5 downto 0) := (others => '0');
begin
	 if rst = '1' then
	 	 count := (others => '0');
	 elsif clk'event and clk = '1' then
	 	 if count = 63 then
	 	 	 count := (others => '0');
	 	 else
	 	 	 count := count+1;
	 	 end if;
	 end if;
	 Counter_out <= count;
end process;
end architecture;

--------------------------------------------------------------------------------
--                          InputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2008)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity InputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(31 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of InputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal expInfty : std_logic := '0';
signal fracZero : std_logic := '0';
signal reprSubNormal : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal infinity : std_logic := '0';
signal zero : std_logic := '0';
signal NaN : std_logic := '0';
signal exnR : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   sX  <= X(31);
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   expInfty  <= '1' when expX = (7 downto 0 => '1') else '0';
   fracZero <= '1' when fracX = (22 downto 0 => '0') else '0';
   reprSubNormal <= fracX(22);
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= fracX(21 downto 0) & '0' when (expZero='1' and reprSubNormal='1')    else fracX;
   fracR <= sfracX;
   -- copy exponent. This will be OK even for subnormals, zero and infty since in such cases the exn bits will prevail
   expR <= expX;
   infinity <= expInfty and fracZero;
   zero <= expZero and not reprSubNormal;
   NaN <= expInfty and not fracZero;
   exnR <= 
           "00" when zero='1' 
      else "10" when infinity='1' 
      else "11" when NaN='1' 
      else "01" ;  -- normal number
   R <= exnR & sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--                         OutputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. Ferrandi  (2009-2012)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity OutputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of OutputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal exnX : std_logic_vector(1 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   exnX  <= X(33 downto 32);
   sX  <= X(31) when (exnX = "01" or exnX = "10" or exnX = "00") else '0';
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= 
      (22 downto 0 => '0') when (exnX = "00") else
      '1' & fracX(22 downto 1) when (expZero = '1' and exnX = "01") else
      fracX when (exnX = "01") else 
      (22 downto 1 => '0') & exnX(0);
   fracR <= sfracX;
   expR <=  
      (7 downto 0 => '0') when (exnX = "00") else
      expX when (exnX = "01") else 
      (7 downto 0 => '1');
   R <= sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_7_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_7_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(2 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_7_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000",
         iS_1 when "001",
         iS_2 when "010",
         iS_3 when "011",
         iS_4 when "100",
         iS_5 when "101",
         iS_6 when "110",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      Y <= s0;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid2599194_RightShifter
--                (RightShifter_24_by_max_26_F250_uid2599196)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid2599194_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid2599194_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_27_f250_uid2599199
--                  (IntAdderAlternative_27_f250_uid2599203)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid2599199 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid2599199 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--              LZCShifter_28_to_28_counting_32_F250_uid2599206
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid2599206 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid2599206 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_34_f250_uid2599209
--                   (IntAdderClassical_34_f250_uid2599211)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid2599209 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid2599209 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                           FPAdd_8_23_uid2599194
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid2599194 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid2599194 is
   component FPAdd_8_23_uid2599194_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid2599199 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid2599206 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid2599209 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid2599194_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid2599199  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid2599206  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid2599209  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   component FPAdd_8_23_uid2599194 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= Y;
   FPAddSubOp_instance: FPAdd_8_23_uid2599194  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_64_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_64_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iS_13 : in std_logic_vector(33 downto 0);
          iS_14 : in std_logic_vector(33 downto 0);
          iS_15 : in std_logic_vector(33 downto 0);
          iS_16 : in std_logic_vector(33 downto 0);
          iS_17 : in std_logic_vector(33 downto 0);
          iS_18 : in std_logic_vector(33 downto 0);
          iS_19 : in std_logic_vector(33 downto 0);
          iS_20 : in std_logic_vector(33 downto 0);
          iS_21 : in std_logic_vector(33 downto 0);
          iS_22 : in std_logic_vector(33 downto 0);
          iS_23 : in std_logic_vector(33 downto 0);
          iS_24 : in std_logic_vector(33 downto 0);
          iS_25 : in std_logic_vector(33 downto 0);
          iS_26 : in std_logic_vector(33 downto 0);
          iS_27 : in std_logic_vector(33 downto 0);
          iS_28 : in std_logic_vector(33 downto 0);
          iS_29 : in std_logic_vector(33 downto 0);
          iS_30 : in std_logic_vector(33 downto 0);
          iS_31 : in std_logic_vector(33 downto 0);
          iS_32 : in std_logic_vector(33 downto 0);
          iS_33 : in std_logic_vector(33 downto 0);
          iS_34 : in std_logic_vector(33 downto 0);
          iS_35 : in std_logic_vector(33 downto 0);
          iS_36 : in std_logic_vector(33 downto 0);
          iS_37 : in std_logic_vector(33 downto 0);
          iS_38 : in std_logic_vector(33 downto 0);
          iS_39 : in std_logic_vector(33 downto 0);
          iS_40 : in std_logic_vector(33 downto 0);
          iS_41 : in std_logic_vector(33 downto 0);
          iS_42 : in std_logic_vector(33 downto 0);
          iS_43 : in std_logic_vector(33 downto 0);
          iS_44 : in std_logic_vector(33 downto 0);
          iS_45 : in std_logic_vector(33 downto 0);
          iS_46 : in std_logic_vector(33 downto 0);
          iS_47 : in std_logic_vector(33 downto 0);
          iS_48 : in std_logic_vector(33 downto 0);
          iS_49 : in std_logic_vector(33 downto 0);
          iS_50 : in std_logic_vector(33 downto 0);
          iS_51 : in std_logic_vector(33 downto 0);
          iS_52 : in std_logic_vector(33 downto 0);
          iS_53 : in std_logic_vector(33 downto 0);
          iS_54 : in std_logic_vector(33 downto 0);
          iS_55 : in std_logic_vector(33 downto 0);
          iS_56 : in std_logic_vector(33 downto 0);
          iS_57 : in std_logic_vector(33 downto 0);
          iS_58 : in std_logic_vector(33 downto 0);
          iS_59 : in std_logic_vector(33 downto 0);
          iS_60 : in std_logic_vector(33 downto 0);
          iS_61 : in std_logic_vector(33 downto 0);
          iS_62 : in std_logic_vector(33 downto 0);
          iS_63 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(5 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_64_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000000",
         iS_1 when "000001",
         iS_2 when "000010",
         iS_3 when "000011",
         iS_4 when "000100",
         iS_5 when "000101",
         iS_6 when "000110",
         iS_7 when "000111",
         iS_8 when "001000",
         iS_9 when "001001",
         iS_10 when "001010",
         iS_11 when "001011",
         iS_12 when "001100",
         iS_13 when "001101",
         iS_14 when "001110",
         iS_15 when "001111",
         iS_16 when "010000",
         iS_17 when "010001",
         iS_18 when "010010",
         iS_19 when "010011",
         iS_20 when "010100",
         iS_21 when "010101",
         iS_22 when "010110",
         iS_23 when "010111",
         iS_24 when "011000",
         iS_25 when "011001",
         iS_26 when "011010",
         iS_27 when "011011",
         iS_28 when "011100",
         iS_29 when "011101",
         iS_30 when "011110",
         iS_31 when "011111",
         iS_32 when "100000",
         iS_33 when "100001",
         iS_34 when "100010",
         iS_35 when "100011",
         iS_36 when "100100",
         iS_37 when "100101",
         iS_38 when "100110",
         iS_39 when "100111",
         iS_40 when "101000",
         iS_41 when "101001",
         iS_42 when "101010",
         iS_43 when "101011",
         iS_44 when "101100",
         iS_45 when "101101",
         iS_46 when "101110",
         iS_47 when "101111",
         iS_48 when "110000",
         iS_49 when "110001",
         iS_50 when "110010",
         iS_51 when "110011",
         iS_52 when "110100",
         iS_53 when "110101",
         iS_54 when "110110",
         iS_55 when "110111",
         iS_56 when "111000",
         iS_57 when "111001",
         iS_58 when "111010",
         iS_59 when "111011",
         iS_60 when "111100",
         iS_61 when "111101",
         iS_62 when "111110",
         iS_63 when "111111",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_63_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_63_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iS_13 : in std_logic_vector(33 downto 0);
          iS_14 : in std_logic_vector(33 downto 0);
          iS_15 : in std_logic_vector(33 downto 0);
          iS_16 : in std_logic_vector(33 downto 0);
          iS_17 : in std_logic_vector(33 downto 0);
          iS_18 : in std_logic_vector(33 downto 0);
          iS_19 : in std_logic_vector(33 downto 0);
          iS_20 : in std_logic_vector(33 downto 0);
          iS_21 : in std_logic_vector(33 downto 0);
          iS_22 : in std_logic_vector(33 downto 0);
          iS_23 : in std_logic_vector(33 downto 0);
          iS_24 : in std_logic_vector(33 downto 0);
          iS_25 : in std_logic_vector(33 downto 0);
          iS_26 : in std_logic_vector(33 downto 0);
          iS_27 : in std_logic_vector(33 downto 0);
          iS_28 : in std_logic_vector(33 downto 0);
          iS_29 : in std_logic_vector(33 downto 0);
          iS_30 : in std_logic_vector(33 downto 0);
          iS_31 : in std_logic_vector(33 downto 0);
          iS_32 : in std_logic_vector(33 downto 0);
          iS_33 : in std_logic_vector(33 downto 0);
          iS_34 : in std_logic_vector(33 downto 0);
          iS_35 : in std_logic_vector(33 downto 0);
          iS_36 : in std_logic_vector(33 downto 0);
          iS_37 : in std_logic_vector(33 downto 0);
          iS_38 : in std_logic_vector(33 downto 0);
          iS_39 : in std_logic_vector(33 downto 0);
          iS_40 : in std_logic_vector(33 downto 0);
          iS_41 : in std_logic_vector(33 downto 0);
          iS_42 : in std_logic_vector(33 downto 0);
          iS_43 : in std_logic_vector(33 downto 0);
          iS_44 : in std_logic_vector(33 downto 0);
          iS_45 : in std_logic_vector(33 downto 0);
          iS_46 : in std_logic_vector(33 downto 0);
          iS_47 : in std_logic_vector(33 downto 0);
          iS_48 : in std_logic_vector(33 downto 0);
          iS_49 : in std_logic_vector(33 downto 0);
          iS_50 : in std_logic_vector(33 downto 0);
          iS_51 : in std_logic_vector(33 downto 0);
          iS_52 : in std_logic_vector(33 downto 0);
          iS_53 : in std_logic_vector(33 downto 0);
          iS_54 : in std_logic_vector(33 downto 0);
          iS_55 : in std_logic_vector(33 downto 0);
          iS_56 : in std_logic_vector(33 downto 0);
          iS_57 : in std_logic_vector(33 downto 0);
          iS_58 : in std_logic_vector(33 downto 0);
          iS_59 : in std_logic_vector(33 downto 0);
          iS_60 : in std_logic_vector(33 downto 0);
          iS_61 : in std_logic_vector(33 downto 0);
          iS_62 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(5 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_63_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000000",
         iS_1 when "000001",
         iS_2 when "000010",
         iS_3 when "000011",
         iS_4 when "000100",
         iS_5 when "000101",
         iS_6 when "000110",
         iS_7 when "000111",
         iS_8 when "001000",
         iS_9 when "001001",
         iS_10 when "001010",
         iS_11 when "001011",
         iS_12 when "001100",
         iS_13 when "001101",
         iS_14 when "001110",
         iS_15 when "001111",
         iS_16 when "010000",
         iS_17 when "010001",
         iS_18 when "010010",
         iS_19 when "010011",
         iS_20 when "010100",
         iS_21 when "010101",
         iS_22 when "010110",
         iS_23 when "010111",
         iS_24 when "011000",
         iS_25 when "011001",
         iS_26 when "011010",
         iS_27 when "011011",
         iS_28 when "011100",
         iS_29 when "011101",
         iS_30 when "011110",
         iS_31 when "011111",
         iS_32 when "100000",
         iS_33 when "100001",
         iS_34 when "100010",
         iS_35 when "100011",
         iS_36 when "100100",
         iS_37 when "100101",
         iS_38 when "100110",
         iS_39 when "100111",
         iS_40 when "101000",
         iS_41 when "101001",
         iS_42 when "101010",
         iS_43 when "101011",
         iS_44 when "101100",
         iS_45 when "101101",
         iS_46 when "101110",
         iS_47 when "101111",
         iS_48 when "110000",
         iS_49 when "110001",
         iS_50 when "110010",
         iS_51 when "110011",
         iS_52 when "110100",
         iS_53 when "110101",
         iS_54 when "110110",
         iS_55 when "110111",
         iS_56 when "111000",
         iS_57 when "111001",
         iS_58 when "111010",
         iS_59 when "111011",
         iS_60 when "111100",
         iS_61 when "111101",
         iS_62 when "111110",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_48_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_48_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iS_13 : in std_logic_vector(33 downto 0);
          iS_14 : in std_logic_vector(33 downto 0);
          iS_15 : in std_logic_vector(33 downto 0);
          iS_16 : in std_logic_vector(33 downto 0);
          iS_17 : in std_logic_vector(33 downto 0);
          iS_18 : in std_logic_vector(33 downto 0);
          iS_19 : in std_logic_vector(33 downto 0);
          iS_20 : in std_logic_vector(33 downto 0);
          iS_21 : in std_logic_vector(33 downto 0);
          iS_22 : in std_logic_vector(33 downto 0);
          iS_23 : in std_logic_vector(33 downto 0);
          iS_24 : in std_logic_vector(33 downto 0);
          iS_25 : in std_logic_vector(33 downto 0);
          iS_26 : in std_logic_vector(33 downto 0);
          iS_27 : in std_logic_vector(33 downto 0);
          iS_28 : in std_logic_vector(33 downto 0);
          iS_29 : in std_logic_vector(33 downto 0);
          iS_30 : in std_logic_vector(33 downto 0);
          iS_31 : in std_logic_vector(33 downto 0);
          iS_32 : in std_logic_vector(33 downto 0);
          iS_33 : in std_logic_vector(33 downto 0);
          iS_34 : in std_logic_vector(33 downto 0);
          iS_35 : in std_logic_vector(33 downto 0);
          iS_36 : in std_logic_vector(33 downto 0);
          iS_37 : in std_logic_vector(33 downto 0);
          iS_38 : in std_logic_vector(33 downto 0);
          iS_39 : in std_logic_vector(33 downto 0);
          iS_40 : in std_logic_vector(33 downto 0);
          iS_41 : in std_logic_vector(33 downto 0);
          iS_42 : in std_logic_vector(33 downto 0);
          iS_43 : in std_logic_vector(33 downto 0);
          iS_44 : in std_logic_vector(33 downto 0);
          iS_45 : in std_logic_vector(33 downto 0);
          iS_46 : in std_logic_vector(33 downto 0);
          iS_47 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(5 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_48_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000000",
         iS_1 when "000001",
         iS_2 when "000010",
         iS_3 when "000011",
         iS_4 when "000100",
         iS_5 when "000101",
         iS_6 when "000110",
         iS_7 when "000111",
         iS_8 when "001000",
         iS_9 when "001001",
         iS_10 when "001010",
         iS_11 when "001011",
         iS_12 when "001100",
         iS_13 when "001101",
         iS_14 when "001110",
         iS_15 when "001111",
         iS_16 when "010000",
         iS_17 when "010001",
         iS_18 when "010010",
         iS_19 when "010011",
         iS_20 when "010100",
         iS_21 when "010101",
         iS_22 when "010110",
         iS_23 when "010111",
         iS_24 when "011000",
         iS_25 when "011001",
         iS_26 when "011010",
         iS_27 when "011011",
         iS_28 when "011100",
         iS_29 when "011101",
         iS_30 when "011110",
         iS_31 when "011111",
         iS_32 when "100000",
         iS_33 when "100001",
         iS_34 when "100010",
         iS_35 when "100011",
         iS_36 when "100100",
         iS_37 when "100101",
         iS_38 when "100110",
         iS_39 when "100111",
         iS_40 when "101000",
         iS_41 when "101001",
         iS_42 when "101010",
         iS_43 when "101011",
         iS_44 when "101100",
         iS_45 when "101101",
         iS_46 when "101110",
         iS_47 when "101111",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_33_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_33_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iS_13 : in std_logic_vector(33 downto 0);
          iS_14 : in std_logic_vector(33 downto 0);
          iS_15 : in std_logic_vector(33 downto 0);
          iS_16 : in std_logic_vector(33 downto 0);
          iS_17 : in std_logic_vector(33 downto 0);
          iS_18 : in std_logic_vector(33 downto 0);
          iS_19 : in std_logic_vector(33 downto 0);
          iS_20 : in std_logic_vector(33 downto 0);
          iS_21 : in std_logic_vector(33 downto 0);
          iS_22 : in std_logic_vector(33 downto 0);
          iS_23 : in std_logic_vector(33 downto 0);
          iS_24 : in std_logic_vector(33 downto 0);
          iS_25 : in std_logic_vector(33 downto 0);
          iS_26 : in std_logic_vector(33 downto 0);
          iS_27 : in std_logic_vector(33 downto 0);
          iS_28 : in std_logic_vector(33 downto 0);
          iS_29 : in std_logic_vector(33 downto 0);
          iS_30 : in std_logic_vector(33 downto 0);
          iS_31 : in std_logic_vector(33 downto 0);
          iS_32 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(5 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_33_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000000",
         iS_1 when "000001",
         iS_2 when "000010",
         iS_3 when "000011",
         iS_4 when "000100",
         iS_5 when "000101",
         iS_6 when "000110",
         iS_7 when "000111",
         iS_8 when "001000",
         iS_9 when "001001",
         iS_10 when "001010",
         iS_11 when "001011",
         iS_12 when "001100",
         iS_13 when "001101",
         iS_14 when "001110",
         iS_15 when "001111",
         iS_16 when "010000",
         iS_17 when "010001",
         iS_18 when "010010",
         iS_19 when "010011",
         iS_20 when "010100",
         iS_21 when "010101",
         iS_22 when "010110",
         iS_23 when "010111",
         iS_24 when "011000",
         iS_25 when "011001",
         iS_26 when "011010",
         iS_27 when "011011",
         iS_28 when "011100",
         iS_29 when "011101",
         iS_30 when "011110",
         iS_31 when "011111",
         iS_32 when "100000",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--          IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid2599624
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid2599624 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          Y : in std_logic_vector(23 downto 0);
          R : out std_logic_vector(47 downto 0)   );
end entity;

architecture arch of IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid2599624 is
signal XX_m2599625 : std_logic_vector(23 downto 0) := (others => '0');
signal YY_m2599625 : std_logic_vector(23 downto 0) := (others => '0');
signal XX : unsigned(-1+24 downto 0) := (others => '0');
signal YY : unsigned(-1+24 downto 0) := (others => '0');
signal RR : unsigned(-1+48 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   XX_m2599625 <= X ;
   YY_m2599625 <= Y ;
   XX <= unsigned(X);
   YY <= unsigned(Y);
   RR <= XX*YY;
   R <= std_logic_vector(RR(47 downto 0));
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_33_f500_uid2599628
--                   (IntAdderClassical_33_f500_uid2599630)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_33_f500_uid2599628 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(32 downto 0);
          Y : in std_logic_vector(32 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(32 downto 0)   );
end entity;

architecture arch of IntAdder_33_f500_uid2599628 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--         FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin 2008-2011
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   component IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid2599624 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             Y : in std_logic_vector(23 downto 0);
             R : out std_logic_vector(47 downto 0)   );
   end component;

   component IntAdder_33_f500_uid2599628 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(32 downto 0);
             Y : in std_logic_vector(32 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(32 downto 0)   );
   end component;

signal sign, sign_d1, sign_d2 : std_logic := '0';
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal expY : std_logic_vector(7 downto 0) := (others => '0');
signal expSumPreSub, expSumPreSub_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal bias, bias_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal expSum : std_logic_vector(9 downto 0) := (others => '0');
signal sigX : std_logic_vector(23 downto 0) := (others => '0');
signal sigY : std_logic_vector(23 downto 0) := (others => '0');
signal sigProd, sigProd_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal excSel : std_logic_vector(3 downto 0) := (others => '0');
signal exc, exc_d1, exc_d2 : std_logic_vector(1 downto 0) := (others => '0');
signal norm : std_logic := '0';
signal expPostNorm : std_logic_vector(9 downto 0) := (others => '0');
signal sigProdExt, sigProdExt_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal expSig, expSig_d1 : std_logic_vector(32 downto 0) := (others => '0');
signal sticky, sticky_d1 : std_logic := '0';
signal guard, guard_d1 : std_logic := '0';
signal round : std_logic := '0';
signal expSigPostRound : std_logic_vector(32 downto 0) := (others => '0');
signal excPostNorm : std_logic_vector(1 downto 0) := (others => '0');
signal finalExc : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            sign_d1 <=  sign;
            sign_d2 <=  sign_d1;
            expSumPreSub_d1 <=  expSumPreSub;
            bias_d1 <=  bias;
            sigProd_d1 <=  sigProd;
            exc_d1 <=  exc;
            exc_d2 <=  exc_d1;
            sigProdExt_d1 <=  sigProdExt;
            expSig_d1 <=  expSig;
            sticky_d1 <=  sticky;
            guard_d1 <=  guard;
         end if;
      end process;
   sign <= X(31) xor Y(31);
   expX <= X(30 downto 23);
   expY <= Y(30 downto 23);
   expSumPreSub <= ("00" & expX) + ("00" & expY);
   bias <= CONV_STD_LOGIC_VECTOR(127,10);
   ----------------Synchro barrier, entering cycle 1----------------
   expSum <= expSumPreSub_d1 - bias_d1;
   ----------------Synchro barrier, entering cycle 0----------------
   sigX <= "1" & X(22 downto 0);
   sigY <= "1" & Y(22 downto 0);
   SignificandMultiplication: IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid2599624  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => sigProd,
                 X => sigX,
                 Y => sigY);
   ----------------Synchro barrier, entering cycle 0----------------
   excSel <= X(33 downto 32) & Y(33 downto 32);
   with excSel select 
   exc <= "00" when  "0000" | "0001" | "0100", 
          "01" when "0101",
          "10" when "0110" | "1001" | "1010" ,
          "11" when others;
   norm <= sigProd_d1(47);
   -- exponent update
   expPostNorm <= expSum + ("000000000" & norm);
   -- significand normalization shift
   sigProdExt <= sigProd_d1(46 downto 0) & "0" when norm='1' else
                         sigProd_d1(45 downto 0) & "00";
   expSig <= expPostNorm & sigProdExt(47 downto 25);
   sticky <= sigProdExt(24);
   guard <= '0' when sigProdExt(23 downto 0)="000000000000000000000000" else '1';
   ----------------Synchro barrier, entering cycle 2----------------
   round <= sticky_d1 and ( (guard_d1 and not(sigProdExt_d1(25))) or (sigProdExt_d1(25) ))  ;
      RoundingAdder: IntAdder_33_f500_uid2599628  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => round,
                 R => expSigPostRound,
                 X => expSig_d1,
                 Y => "000000000000000000000000000000000");
   with expSigPostRound(32 downto 31) select
   excPostNorm <=  "01"  when  "00",
                               "10"             when "01", 
                               "00"             when "11"|"10",
                               "11"             when others;
   with exc_d2 select 
   finalExc <= exc_d2 when  "11"|"10"|"00",
                       excPostNorm when others; 
   R <= finalExc & sign_d2 & expSigPostRound(30 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid2599931_RightShifter
--                (RightShifter_24_by_max_26_F250_uid2599933)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid2599931_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid2599931_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_27_f250_uid2599936
--                  (IntAdderAlternative_27_f250_uid2599940)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid2599936 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid2599936 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--              LZCShifter_28_to_28_counting_32_F250_uid2599943
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid2599943 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid2599943 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_34_f250_uid2599946
--                   (IntAdderClassical_34_f250_uid2599948)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid2599946 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid2599946 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                           FPAdd_8_23_uid2599931
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid2599931 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid2599931 is
   component FPAdd_8_23_uid2599931_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid2599936 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid2599943 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid2599946 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid2599931_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid2599936  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid2599943  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid2599946  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
   component FPAdd_8_23_uid2599931 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= (Y(Y'length-1 downto Y'length-2)) & (not Y(Y'length-3)) & Y(Y'length-4 downto 0);
   FPAddSubOp_instance: FPAdd_8_23_uid2599931  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_47_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_47_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iS_13 : in std_logic_vector(33 downto 0);
          iS_14 : in std_logic_vector(33 downto 0);
          iS_15 : in std_logic_vector(33 downto 0);
          iS_16 : in std_logic_vector(33 downto 0);
          iS_17 : in std_logic_vector(33 downto 0);
          iS_18 : in std_logic_vector(33 downto 0);
          iS_19 : in std_logic_vector(33 downto 0);
          iS_20 : in std_logic_vector(33 downto 0);
          iS_21 : in std_logic_vector(33 downto 0);
          iS_22 : in std_logic_vector(33 downto 0);
          iS_23 : in std_logic_vector(33 downto 0);
          iS_24 : in std_logic_vector(33 downto 0);
          iS_25 : in std_logic_vector(33 downto 0);
          iS_26 : in std_logic_vector(33 downto 0);
          iS_27 : in std_logic_vector(33 downto 0);
          iS_28 : in std_logic_vector(33 downto 0);
          iS_29 : in std_logic_vector(33 downto 0);
          iS_30 : in std_logic_vector(33 downto 0);
          iS_31 : in std_logic_vector(33 downto 0);
          iS_32 : in std_logic_vector(33 downto 0);
          iS_33 : in std_logic_vector(33 downto 0);
          iS_34 : in std_logic_vector(33 downto 0);
          iS_35 : in std_logic_vector(33 downto 0);
          iS_36 : in std_logic_vector(33 downto 0);
          iS_37 : in std_logic_vector(33 downto 0);
          iS_38 : in std_logic_vector(33 downto 0);
          iS_39 : in std_logic_vector(33 downto 0);
          iS_40 : in std_logic_vector(33 downto 0);
          iS_41 : in std_logic_vector(33 downto 0);
          iS_42 : in std_logic_vector(33 downto 0);
          iS_43 : in std_logic_vector(33 downto 0);
          iS_44 : in std_logic_vector(33 downto 0);
          iS_45 : in std_logic_vector(33 downto 0);
          iS_46 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(5 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_47_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000000",
         iS_1 when "000001",
         iS_2 when "000010",
         iS_3 when "000011",
         iS_4 when "000100",
         iS_5 when "000101",
         iS_6 when "000110",
         iS_7 when "000111",
         iS_8 when "001000",
         iS_9 when "001001",
         iS_10 when "001010",
         iS_11 when "001011",
         iS_12 when "001100",
         iS_13 when "001101",
         iS_14 when "001110",
         iS_15 when "001111",
         iS_16 when "010000",
         iS_17 when "010001",
         iS_18 when "010010",
         iS_19 when "010011",
         iS_20 when "010100",
         iS_21 when "010101",
         iS_22 when "010110",
         iS_23 when "010111",
         iS_24 when "011000",
         iS_25 when "011001",
         iS_26 when "011010",
         iS_27 when "011011",
         iS_28 when "011100",
         iS_29 when "011101",
         iS_30 when "011110",
         iS_31 when "011111",
         iS_32 when "100000",
         iS_33 when "100001",
         iS_34 when "100010",
         iS_35 when "100011",
         iS_36 when "100100",
         iS_37 when "100101",
         iS_38 when "100110",
         iS_39 when "100111",
         iS_40 when "101000",
         iS_41 when "101001",
         iS_42 when "101010",
         iS_43 when "101011",
         iS_44 when "101100",
         iS_45 when "101101",
         iS_46 when "101110",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_34_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_34_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iS_13 : in std_logic_vector(33 downto 0);
          iS_14 : in std_logic_vector(33 downto 0);
          iS_15 : in std_logic_vector(33 downto 0);
          iS_16 : in std_logic_vector(33 downto 0);
          iS_17 : in std_logic_vector(33 downto 0);
          iS_18 : in std_logic_vector(33 downto 0);
          iS_19 : in std_logic_vector(33 downto 0);
          iS_20 : in std_logic_vector(33 downto 0);
          iS_21 : in std_logic_vector(33 downto 0);
          iS_22 : in std_logic_vector(33 downto 0);
          iS_23 : in std_logic_vector(33 downto 0);
          iS_24 : in std_logic_vector(33 downto 0);
          iS_25 : in std_logic_vector(33 downto 0);
          iS_26 : in std_logic_vector(33 downto 0);
          iS_27 : in std_logic_vector(33 downto 0);
          iS_28 : in std_logic_vector(33 downto 0);
          iS_29 : in std_logic_vector(33 downto 0);
          iS_30 : in std_logic_vector(33 downto 0);
          iS_31 : in std_logic_vector(33 downto 0);
          iS_32 : in std_logic_vector(33 downto 0);
          iS_33 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(5 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_34_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000000",
         iS_1 when "000001",
         iS_2 when "000010",
         iS_3 when "000011",
         iS_4 when "000100",
         iS_5 when "000101",
         iS_6 when "000110",
         iS_7 when "000111",
         iS_8 when "001000",
         iS_9 when "001001",
         iS_10 when "001010",
         iS_11 when "001011",
         iS_12 when "001100",
         iS_13 when "001101",
         iS_14 when "001110",
         iS_15 when "001111",
         iS_16 when "010000",
         iS_17 when "010001",
         iS_18 when "010010",
         iS_19 when "010011",
         iS_20 when "010100",
         iS_21 when "010101",
         iS_22 when "010110",
         iS_23 when "010111",
         iS_24 when "011000",
         iS_25 when "011001",
         iS_26 when "011010",
         iS_27 when "011011",
         iS_28 when "011100",
         iS_29 when "011101",
         iS_30 when "011110",
         iS_31 when "011111",
         iS_32 when "100000",
         iS_33 when "100001",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--                      Constant_float_8_23_1_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_1_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_1_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111100000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                      Constant_float_8_23_0_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_0_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_0_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0000000000000000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_cosnpi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosnpi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosnpi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_sinnpi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinnpi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinnpi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn3_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn3_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn3_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn3_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn3_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn3_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_cosnpi_div_2_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosnpi_div_2_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosnpi_div_2_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0000000000000000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_sinnpi_div_2_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinnpi_div_2_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinnpi_div_2_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111100000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn5_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn5_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn5_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn5_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn5_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn5_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn3_mult_pi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn3_mult_pi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn3_mult_pi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn3_mult_pi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn3_mult_pi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn3_mult_pi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn7_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn7_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn7_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn7_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn7_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn7_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_cosnpi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosnpi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosnpi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_sinnpi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinnpi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinnpi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 19 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      Y <= s18;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 14 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      Y <= s13;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      Y <= s1;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "101" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "110" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "001" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "010" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "011" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when "111000",
      "000" when "111001",
      "000" when "111010",
      "000" when "111011",
      "000" when "111100",
      "000" when "111101",
      "100" when "111110",
      "000" when "111111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "101" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "110" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "001" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "010" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "011" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when "111000",
      "000" when "111001",
      "000" when "111010",
      "000" when "111011",
      "000" when "111100",
      "000" when "111101",
      "100" when "111110",
      "000" when "111111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "010" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "011" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "100" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "101" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "110" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when "111000",
      "001" when "111001",
      "000" when "111010",
      "000" when "111011",
      "000" when "111100",
      "000" when "111101",
      "000" when "111110",
      "000" when "111111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "010" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "011" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "100" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "101" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "110" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when "111000",
      "001" when "111001",
      "000" when "111010",
      "000" when "111011",
      "000" when "111100",
      "000" when "111101",
      "000" when "111110",
      "000" when "111111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "100" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "101" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "110" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "001" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "010" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "011" when "111000",
      "000" when "111001",
      "000" when "111010",
      "000" when "111011",
      "000" when "111100",
      "000" when "111101",
      "000" when "111110",
      "000" when "111111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "100" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "101" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "110" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "001" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "010" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "011" when "111000",
      "000" when "111001",
      "000" when "111010",
      "000" when "111011",
      "000" when "111100",
      "000" when "111101",
      "000" when "111110",
      "000" when "111111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "010" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "011" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "100" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "101" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "110" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when "111000",
      "000" when "111001",
      "000" when "111010",
      "000" when "111011",
      "000" when "111100",
      "001" when "111101",
      "000" when "111110",
      "000" when "111111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "010" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "011" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "100" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "101" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "110" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when "111000",
      "000" when "111001",
      "000" when "111010",
      "000" when "111011",
      "000" when "111100",
      "000" when "111101",
      "001" when "111110",
      "000" when "111111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "101" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "110" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "001" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "010" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "011" when "110110",
      "000" when "110111",
      "000" when "111000",
      "000" when "111001",
      "000" when "111010",
      "000" when "111011",
      "000" when "111100",
      "000" when "111101",
      "000" when "111110",
      "100" when "111111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "101" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "110" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "001" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "010" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "011" when "110110",
      "000" when "110111",
      "000" when "111000",
      "000" when "111001",
      "000" when "111010",
      "000" when "111011",
      "000" when "111100",
      "000" when "111101",
      "000" when "111110",
      "100" when "111111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "010" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "011" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "100" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "101" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "110" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when "111000",
      "000" when "111001",
      "001" when "111010",
      "000" when "111011",
      "000" when "111100",
      "000" when "111101",
      "000" when "111110",
      "000" when "111111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "010" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "011" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "100" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "101" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "110" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when "111000",
      "000" when "111001",
      "000" when "111010",
      "001" when "111011",
      "000" when "111100",
      "000" when "111101",
      "000" when "111110",
      "000" when "111111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "100" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "101" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "110" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "001" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "010" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when "111000",
      "011" when "111001",
      "000" when "111010",
      "000" when "111011",
      "000" when "111100",
      "000" when "111101",
      "000" when "111110",
      "000" when "111111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "100" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "101" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "110" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "001" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "010" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when "111000",
      "000" when "111001",
      "011" when "111010",
      "000" when "111011",
      "000" when "111100",
      "000" when "111101",
      "000" when "111110",
      "000" when "111111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "010" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "011" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "100" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "101" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "110" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when "111000",
      "000" when "111001",
      "000" when "111010",
      "000" when "111011",
      "000" when "111100",
      "000" when "111101",
      "001" when "111110",
      "000" when "111111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "010" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "011" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "100" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "101" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "110" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when "111000",
      "000" when "111001",
      "000" when "111010",
      "000" when "111011",
      "000" when "111100",
      "000" when "111101",
      "000" when "111110",
      "001" when "111111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "101" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "110" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "001" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "010" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "011" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when "111000",
      "000" when "111001",
      "000" when "111010",
      "000" when "111011",
      "000" when "111100",
      "000" when "111101",
      "100" when "111110",
      "000" when "111111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "101" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "110" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "001" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "010" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "011" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when "111000",
      "000" when "111001",
      "000" when "111010",
      "000" when "111011",
      "000" when "111100",
      "000" when "111101",
      "100" when "111110",
      "000" when "111111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "010" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "011" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "100" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "101" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "110" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when "111000",
      "001" when "111001",
      "000" when "111010",
      "000" when "111011",
      "000" when "111100",
      "000" when "111101",
      "000" when "111110",
      "000" when "111111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "010" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "011" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "100" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "101" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "110" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when "111000",
      "000" when "111001",
      "001" when "111010",
      "000" when "111011",
      "000" when "111100",
      "000" when "111101",
      "000" when "111110",
      "000" when "111111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "100" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "101" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "110" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "001" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "010" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when "111000",
      "011" when "111001",
      "000" when "111010",
      "000" when "111011",
      "000" when "111100",
      "000" when "111101",
      "000" when "111110",
      "000" when "111111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "100" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "101" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "110" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "001" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "010" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "011" when "111000",
      "000" when "111001",
      "000" when "111010",
      "000" when "111011",
      "000" when "111100",
      "000" when "111101",
      "000" when "111110",
      "000" when "111111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "010" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "011" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "100" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "101" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "110" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when "111000",
      "000" when "111001",
      "000" when "111010",
      "000" when "111011",
      "001" when "111100",
      "000" when "111101",
      "000" when "111110",
      "000" when "111111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "010" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "011" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "100" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "101" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "110" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when "111000",
      "000" when "111001",
      "000" when "111010",
      "000" when "111011",
      "000" when "111100",
      "000" when "111101",
      "001" when "111110",
      "000" when "111111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "101" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "110" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "001" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "010" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "011" when "110110",
      "000" when "110111",
      "000" when "111000",
      "000" when "111001",
      "000" when "111010",
      "000" when "111011",
      "000" when "111100",
      "000" when "111101",
      "000" when "111110",
      "100" when "111111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "101" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "110" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "001" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "010" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "011" when "110110",
      "000" when "110111",
      "000" when "111000",
      "000" when "111001",
      "000" when "111010",
      "000" when "111011",
      "000" when "111100",
      "000" when "111101",
      "000" when "111110",
      "100" when "111111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "010" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "011" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "100" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "101" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "110" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when "111000",
      "000" when "111001",
      "000" when "111010",
      "001" when "111011",
      "000" when "111100",
      "000" when "111101",
      "000" when "111110",
      "000" when "111111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "010" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "011" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "100" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "101" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "110" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when "111000",
      "000" when "111001",
      "000" when "111010",
      "000" when "111011",
      "001" when "111100",
      "000" when "111101",
      "000" when "111110",
      "000" when "111111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "100" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "101" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "110" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "001" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "010" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when "111000",
      "000" when "111001",
      "000" when "111010",
      "011" when "111011",
      "000" when "111100",
      "000" when "111101",
      "000" when "111110",
      "000" when "111111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "101" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "110" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "001" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "010" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "011" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when "111000",
      "000" when "111001",
      "000" when "111010",
      "100" when "111011",
      "000" when "111100",
      "000" when "111101",
      "000" when "111110",
      "000" when "111111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "010" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "011" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "100" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "101" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "110" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when "111000",
      "000" when "111001",
      "000" when "111010",
      "000" when "111011",
      "000" when "111100",
      "000" when "111101",
      "001" when "111110",
      "000" when "111111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "010" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "011" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "100" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "101" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "110" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when "111000",
      "000" when "111001",
      "000" when "111010",
      "000" when "111011",
      "000" when "111100",
      "000" when "111101",
      "000" when "111110",
      "001" when "111111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Add2_5_impl_0_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add2_5_impl_0_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add2_5_impl_0_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "010000" when "000000",
      "011110" when "000001",
      "010110" when "000010",
      "011000" when "000011",
      "100001" when "000100",
      "100010" when "000101",
      "001111" when "000110",
      "111110" when "000111",
      "101011" when "001000",
      "100100" when "001001",
      "111011" when "001010",
      "001010" when "001011",
      "100111" when "001100",
      "110010" when "001101",
      "001100" when "001110",
      "001101" when "001111",
      "001011" when "010000",
      "101001" when "010001",
      "101111" when "010010",
      "110110" when "010011",
      "110001" when "010100",
      "001110" when "010101",
      "111100" when "010110",
      "011010" when "010111",
      "101110" when "011000",
      "010011" when "011001",
      "100101" when "011010",
      "010101" when "011011",
      "100110" when "011100",
      "111001" when "011101",
      "011100" when "011110",
      "000000" when "011111",
      "100011" when "100000",
      "011001" when "100001",
      "011011" when "100010",
      "110100" when "100011",
      "110011" when "100100",
      "100000" when "100101",
      "011111" when "100110",
      "110101" when "100111",
      "011101" when "101000",
      "010001" when "101001",
      "010111" when "101010",
      "110000" when "101011",
      "110111" when "101100",
      "111010" when "101101",
      "000000" when "101110",
      "000001" when "101111",
      "001000" when "110000",
      "010010" when "110001",
      "010100" when "110010",
      "000101" when "110011",
      "000100" when "110100",
      "000110" when "110101",
      "111000" when "110110",
      "101101" when "110111",
      "101100" when "111000",
      "000010" when "111001",
      "001001" when "111010",
      "000111" when "111011",
      "111101" when "111100",
      "101000" when "111101",
      "101010" when "111110",
      "000011" when "111111",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Add2_5_impl_0_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add2_5_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add2_5_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Add2_5_impl_0_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Add2_5_impl_0_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Add2_5_impl_1_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add2_5_impl_1_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add2_5_impl_1_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "001100" when "000000",
      "010011" when "000001",
      "011101" when "000010",
      "011110" when "000011",
      "010010" when "000100",
      "100011" when "000101",
      "001010" when "000110",
      "111100" when "000111",
      "100101" when "001000",
      "011100" when "001001",
      "111001" when "001010",
      "010001" when "001011",
      "100001" when "001100",
      "101111" when "001101",
      "101110" when "001110",
      "111000" when "001111",
      "101100" when "010000",
      "100110" when "010001",
      "101000" when "010010",
      "110010" when "010011",
      "101101" when "010100",
      "001011" when "010101",
      "111011" when "010110",
      "010000" when "010111",
      "101001" when "011000",
      "001110" when "011001",
      "111101" when "011010",
      "111010" when "011011",
      "100000" when "011100",
      "110100" when "011101",
      "010111" when "011110",
      "000000" when "011111",
      "011010" when "100000",
      "011111" when "100001",
      "010101" when "100010",
      "110001" when "100011",
      "110000" when "100100",
      "011011" when "100101",
      "011001" when "100110",
      "110011" when "100111",
      "011000" when "101000",
      "001101" when "101001",
      "001111" when "101010",
      "101011" when "101011",
      "110101" when "101100",
      "110111" when "101101",
      "000000" when "101110",
      "000001" when "101111",
      "001000" when "110000",
      "010100" when "110001",
      "010110" when "110010",
      "000101" when "110011",
      "000100" when "110100",
      "000110" when "110101",
      "110110" when "110110",
      "100111" when "110111",
      "101010" when "111000",
      "000010" when "111001",
      "001001" when "111010",
      "000111" when "111011",
      "111110" when "111100",
      "100010" when "111101",
      "100100" when "111110",
      "000011" when "111111",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Add2_5_impl_1_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add2_5_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add2_5_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Add2_5_impl_1_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Add2_5_impl_1_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Add2_6_impl_0_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add2_6_impl_0_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add2_6_impl_0_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "100011" when "000000",
      "100001" when "000001",
      "100110" when "000010",
      "000000" when "000011",
      "000000" when "000100",
      "011001" when "000101",
      "100111" when "000110",
      "001011" when "000111",
      "000000" when "001000",
      "010010" when "001001",
      "001110" when "001010",
      "011101" when "001011",
      "000000" when "001100",
      "000000" when "001101",
      "011100" when "001110",
      "100010" when "001111",
      "100100" when "010000",
      "101110" when "010001",
      "010000" when "010010",
      "101111" when "010011",
      "101101" when "010100",
      "000000" when "010101",
      "000000" when "010110",
      "101010" when "010111",
      "100000" when "011000",
      "001100" when "011001",
      "001010" when "011010",
      "001111" when "011011",
      "010001" when "011100",
      "101000" when "011101",
      "101011" when "011110",
      "000000" when "011111",
      "010111" when "100000",
      "001101" when "100001",
      "100101" when "100010",
      "010100" when "100011",
      "011111" when "100100",
      "011010" when "100101",
      "101001" when "100110",
      "101100" when "100111",
      "000000" when "101000",
      "000000" when "101001",
      "010011" when "101010",
      "011000" when "101011",
      "011011" when "101100",
      "010110" when "101101",
      "000001" when "101110",
      "000010" when "101111",
      "011110" when "110000",
      "000000" when "110001",
      "000000" when "110010",
      "001000" when "110011",
      "001001" when "110100",
      "000101" when "110101",
      "000000" when "110110",
      "010101" when "110111",
      "000000" when "111000",
      "000011" when "111001",
      "000000" when "111010",
      "000000" when "111011",
      "000100" when "111100",
      "000111" when "111101",
      "000110" when "111110",
      "000000" when "111111",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Add2_6_impl_0_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add2_6_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add2_6_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Add2_6_impl_0_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Add2_6_impl_0_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Add2_6_impl_1_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add2_6_impl_1_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add2_6_impl_1_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "100000" when "000000",
      "011111" when "000001",
      "100011" when "000010",
      "000000" when "000011",
      "000000" when "000100",
      "010110" when "000101",
      "100110" when "000110",
      "001010" when "000111",
      "000000" when "001000",
      "011001" when "001001",
      "001011" when "001010",
      "011010" when "001011",
      "000000" when "001100",
      "000000" when "001101",
      "011100" when "001110",
      "100001" when "001111",
      "100010" when "010000",
      "101111" when "010001",
      "001110" when "010010",
      "001100" when "010011",
      "101101" when "010100",
      "000000" when "010101",
      "000000" when "010110",
      "001101" when "010111",
      "101001" when "011000",
      "101110" when "011001",
      "100101" when "011010",
      "010001" when "011011",
      "010000" when "011100",
      "100111" when "011101",
      "101011" when "011110",
      "000000" when "011111",
      "010101" when "100000",
      "001111" when "100001",
      "100100" when "100010",
      "010010" when "100011",
      "011011" when "100100",
      "101100" when "100101",
      "101010" when "100110",
      "101000" when "100111",
      "000000" when "101000",
      "000000" when "101001",
      "010111" when "101010",
      "011000" when "101011",
      "011110" when "101100",
      "010011" when "101101",
      "000010" when "101110",
      "000011" when "101111",
      "011101" when "110000",
      "000000" when "110001",
      "000000" when "110010",
      "001000" when "110011",
      "001001" when "110100",
      "000101" when "110101",
      "000000" when "110110",
      "010100" when "110111",
      "000001" when "111000",
      "000100" when "111001",
      "000000" when "111010",
      "000000" when "111011",
      "000000" when "111100",
      "000111" when "111101",
      "000110" when "111110",
      "000000" when "111111",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Add2_6_impl_1_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add2_6_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add2_6_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Add2_6_impl_1_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Add2_6_impl_1_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Add11_6_impl_0_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add11_6_impl_0_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add11_6_impl_0_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "011011" when "000000",
      "010111" when "000001",
      "000000" when "000010",
      "000000" when "000011",
      "000000" when "000100",
      "010101" when "000101",
      "011111" when "000110",
      "010110" when "000111",
      "000000" when "001000",
      "100000" when "001001",
      "001000" when "001010",
      "000000" when "001011",
      "000000" when "001100",
      "000000" when "001101",
      "000111" when "001110",
      "010000" when "001111",
      "000110" when "010000",
      "000000" when "010001",
      "000000" when "010010",
      "010010" when "010011",
      "000000" when "010100",
      "000000" when "010101",
      "000000" when "010110",
      "011110" when "010111",
      "000100" when "011000",
      "000101" when "011001",
      "000000" when "011010",
      "000000" when "011011",
      "011001" when "011100",
      "011100" when "011101",
      "000000" when "011110",
      "000000" when "011111",
      "000000" when "100000",
      "001101" when "100001",
      "011000" when "100010",
      "000000" when "100011",
      "000000" when "100100",
      "001011" when "100101",
      "010100" when "100110",
      "000000" when "100111",
      "000000" when "101000",
      "000000" when "101001",
      "010001" when "101010",
      "001100" when "101011",
      "001110" when "101100",
      "000000" when "101101",
      "001010" when "101110",
      "001111" when "101111",
      "000000" when "110000",
      "000000" when "110001",
      "000000" when "110010",
      "010011" when "110011",
      "001001" when "110100",
      "011010" when "110101",
      "000000" when "110110",
      "011101" when "110111",
      "000000" when "111000",
      "000000" when "111001",
      "000000" when "111010",
      "000000" when "111011",
      "000001" when "111100",
      "000010" when "111101",
      "000011" when "111110",
      "000000" when "111111",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Add11_6_impl_0_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add11_6_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add11_6_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Add11_6_impl_0_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Add11_6_impl_0_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Add11_6_impl_1_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add11_6_impl_1_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add11_6_impl_1_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "011011" when "000000",
      "010110" when "000001",
      "000000" when "000010",
      "000000" when "000011",
      "000000" when "000100",
      "010011" when "000101",
      "100000" when "000110",
      "010100" when "000111",
      "000000" when "001000",
      "011111" when "001001",
      "000111" when "001010",
      "000000" when "001011",
      "000000" when "001100",
      "000000" when "001101",
      "000101" when "001110",
      "010101" when "001111",
      "000100" when "010000",
      "000000" when "010001",
      "000000" when "010010",
      "001111" when "010011",
      "000000" when "010100",
      "000000" when "010101",
      "000000" when "010110",
      "000110" when "010111",
      "011010" when "011000",
      "011110" when "011001",
      "000000" when "011010",
      "000000" when "011011",
      "010111" when "011100",
      "011100" when "011101",
      "000000" when "011110",
      "000000" when "011111",
      "000000" when "100000",
      "001011" when "100001",
      "011000" when "100010",
      "000000" when "100011",
      "000000" when "100100",
      "001001" when "100101",
      "010010" when "100110",
      "000000" when "100111",
      "000000" when "101000",
      "000000" when "101001",
      "001101" when "101010",
      "010001" when "101011",
      "001100" when "101100",
      "000000" when "101101",
      "001000" when "101110",
      "001110" when "101111",
      "000000" when "110000",
      "000000" when "110001",
      "000000" when "110010",
      "010000" when "110011",
      "001010" when "110100",
      "011001" when "110101",
      "000000" when "110110",
      "011101" when "110111",
      "000000" when "111000",
      "000000" when "111001",
      "000000" when "111010",
      "000000" when "111011",
      "000001" when "111100",
      "000010" when "111101",
      "000011" when "111110",
      "000000" when "111111",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Add11_6_impl_1_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add11_6_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add11_6_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Add11_6_impl_1_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Add11_6_impl_1_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Subtract2_6_impl_0_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract2_6_impl_0_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract2_6_impl_0_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "100001" when "000000",
      "001011" when "000001",
      "011000" when "000010",
      "011100" when "000011",
      "100100" when "000100",
      "100000" when "000101",
      "100111" when "000110",
      "111011" when "000111",
      "001100" when "001000",
      "101111" when "001001",
      "111101" when "001010",
      "010011" when "001011",
      "100110" when "001100",
      "110000" when "001101",
      "001101" when "001110",
      "010000" when "001111",
      "001110" when "010000",
      "111100" when "010001",
      "111001" when "010010",
      "110011" when "010011",
      "111000" when "010100",
      "010010" when "010101",
      "111110" when "010110",
      "010001" when "010111",
      "101100" when "011000",
      "101010" when "011001",
      "001111" when "011010",
      "110100" when "011011",
      "100101" when "011100",
      "110111" when "011101",
      "110101" when "011110",
      "000000" when "011111",
      "010110" when "100000",
      "011101" when "100001",
      "011110" when "100010",
      "101011" when "100011",
      "011001" when "100100",
      "100011" when "100101",
      "100010" when "100110",
      "110010" when "100111",
      "110110" when "101000",
      "010100" when "101001",
      "011011" when "101010",
      "101110" when "101011",
      "011111" when "101100",
      "110001" when "101101",
      "000001" when "101110",
      "000010" when "101111",
      "001001" when "110000",
      "010101" when "110001",
      "010111" when "110010",
      "000111" when "110011",
      "000101" when "110100",
      "001000" when "110101",
      "101001" when "110110",
      "101101" when "110111",
      "011010" when "111000",
      "000011" when "111001",
      "001010" when "111010",
      "000000" when "111011",
      "111010" when "111100",
      "101000" when "111101",
      "000110" when "111110",
      "000100" when "111111",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Subtract2_6_impl_0_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract2_6_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract2_6_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Subtract2_6_impl_0_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Subtract2_6_impl_0_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Subtract2_6_impl_1_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract2_6_impl_1_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract2_6_impl_1_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "011000" when "000000",
      "010110" when "000001",
      "010010" when "000010",
      "100001" when "000011",
      "010111" when "000100",
      "011100" when "000101",
      "100110" when "000110",
      "111100" when "000111",
      "001011" when "001000",
      "101110" when "001001",
      "001100" when "001010",
      "010000" when "001011",
      "100100" when "001100",
      "101011" when "001101",
      "101111" when "001110",
      "111010" when "001111",
      "110111" when "010000",
      "111101" when "010001",
      "111011" when "010010",
      "110001" when "010011",
      "111001" when "010100",
      "001111" when "010101",
      "001101" when "010110",
      "001110" when "010111",
      "101101" when "011000",
      "101000" when "011001",
      "111000" when "011010",
      "110100" when "011011",
      "011111" when "011100",
      "110011" when "011101",
      "110101" when "011110",
      "000000" when "011111",
      "010100" when "100000",
      "100010" when "100001",
      "100011" when "100010",
      "101001" when "100011",
      "010011" when "100100",
      "011110" when "100101",
      "011101" when "100110",
      "110010" when "100111",
      "110110" when "101000",
      "010001" when "101001",
      "010101" when "101010",
      "101100" when "101011",
      "011010" when "101100",
      "110000" when "101101",
      "000000" when "101110",
      "000001" when "101111",
      "001001" when "110000",
      "011001" when "110001",
      "011011" when "110010",
      "000111" when "110011",
      "000101" when "110100",
      "001000" when "110101",
      "100111" when "110110",
      "101010" when "110111",
      "100000" when "111000",
      "000010" when "111001",
      "001010" when "111010",
      "000011" when "111011",
      "111110" when "111100",
      "100101" when "111101",
      "000110" when "111110",
      "000100" when "111111",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Subtract2_6_impl_1_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract2_6_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract2_6_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Subtract2_6_impl_1_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Subtract2_6_impl_1_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Subtract3_6_impl_0_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract3_6_impl_0_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract3_6_impl_0_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "100001" when "000000",
      "100000" when "000001",
      "010101" when "000010",
      "000000" when "000011",
      "000000" when "000100",
      "010011" when "000101",
      "100101" when "000110",
      "011100" when "000111",
      "000000" when "001000",
      "001101" when "001001",
      "001100" when "001010",
      "001011" when "001011",
      "000000" when "001100",
      "000000" when "001101",
      "001111" when "001110",
      "011011" when "001111",
      "001110" when "010000",
      "000000" when "010001",
      "100010" when "010010",
      "011111" when "010011",
      "101110" when "010100",
      "000000" when "010101",
      "000000" when "010110",
      "101001" when "010111",
      "011110" when "011000",
      "001010" when "011001",
      "000000" when "011010",
      "010010" when "011011",
      "100011" when "011100",
      "100111" when "011101",
      "101011" when "011110",
      "000000" when "011111",
      "010000" when "100000",
      "010111" when "100001",
      "010100" when "100010",
      "000000" when "100011",
      "011010" when "100100",
      "100110" when "100101",
      "010110" when "100110",
      "101100" when "100111",
      "000000" when "101000",
      "000000" when "101001",
      "011101" when "101010",
      "010001" when "101011",
      "011000" when "101100",
      "101101" when "101101",
      "000001" when "101110",
      "000010" when "101111",
      "011001" when "110000",
      "000000" when "110001",
      "000000" when "110010",
      "000110" when "110011",
      "001000" when "110100",
      "100100" when "110101",
      "101010" when "110110",
      "101000" when "110111",
      "000000" when "111000",
      "000011" when "111001",
      "000000" when "111010",
      "000000" when "111011",
      "000100" when "111100",
      "000101" when "111101",
      "001001" when "111110",
      "000111" when "111111",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Subtract3_6_impl_0_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract3_6_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract3_6_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Subtract3_6_impl_0_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Subtract3_6_impl_0_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Subtract3_6_impl_1_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract3_6_impl_1_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract3_6_impl_1_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "011111" when "000000",
      "011100" when "000001",
      "011010" when "000010",
      "000000" when "000011",
      "000000" when "000100",
      "010001" when "000101",
      "100100" when "000110",
      "011101" when "000111",
      "000000" when "001000",
      "001100" when "001001",
      "001010" when "001010",
      "010101" when "001011",
      "000000" when "001100",
      "000000" when "001101",
      "001011" when "001110",
      "011110" when "001111",
      "001101" when "010000",
      "000000" when "010001",
      "100000" when "010010",
      "011001" when "010011",
      "001110" when "010100",
      "000000" when "010101",
      "000000" when "010110",
      "001111" when "010111",
      "101001" when "011000",
      "100001" when "011001",
      "000000" when "011010",
      "101110" when "011011",
      "100010" when "011100",
      "100101" when "011101",
      "101100" when "011110",
      "000000" when "011111",
      "010000" when "100000",
      "010100" when "100001",
      "101101" when "100010",
      "000000" when "100011",
      "010110" when "100100",
      "100110" when "100101",
      "010010" when "100110",
      "101000" when "100111",
      "000000" when "101000",
      "000000" when "101001",
      "011000" when "101010",
      "010011" when "101011",
      "011011" when "101100",
      "101010" when "101101",
      "000010" when "101110",
      "000011" when "101111",
      "010111" when "110000",
      "000000" when "110001",
      "000000" when "110010",
      "000110" when "110011",
      "001000" when "110100",
      "100011" when "110101",
      "101011" when "110110",
      "100111" when "110111",
      "000001" when "111000",
      "000100" when "111001",
      "000000" when "111010",
      "000000" when "111011",
      "000000" when "111100",
      "000101" when "111101",
      "001001" when "111110",
      "000111" when "111111",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Subtract3_6_impl_1_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract3_6_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract3_6_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Subtract3_6_impl_1_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Subtract3_6_impl_1_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--        GenericLut_LUTData_MUX_Subtract12_6_impl_0_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract12_6_impl_0_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract12_6_impl_0_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "010110" when "000000",
      "010111" when "000001",
      "000000" when "000010",
      "000000" when "000011",
      "000000" when "000100",
      "010010" when "000101",
      "100000" when "000110",
      "010101" when "000111",
      "000000" when "001000",
      "000111" when "001001",
      "001110" when "001010",
      "000000" when "001011",
      "000000" when "001100",
      "000000" when "001101",
      "100001" when "001110",
      "001101" when "001111",
      "010011" when "010000",
      "000000" when "010001",
      "010100" when "010010",
      "011001" when "010011",
      "000000" when "010100",
      "000000" when "010101",
      "000000" when "010110",
      "011111" when "010111",
      "000011" when "011000",
      "000100" when "011001",
      "000000" when "011010",
      "000110" when "011011",
      "011110" when "011100",
      "011011" when "011101",
      "000000" when "011110",
      "000000" when "011111",
      "000000" when "100000",
      "000101" when "100001",
      "011000" when "100010",
      "000000" when "100011",
      "011010" when "100100",
      "011100" when "100101",
      "010001" when "100110",
      "000000" when "100111",
      "000000" when "101000",
      "000000" when "101001",
      "001000" when "101010",
      "001100" when "101011",
      "000000" when "101100",
      "001001" when "101101",
      "001010" when "101110",
      "001111" when "101111",
      "000000" when "110000",
      "000000" when "110001",
      "000000" when "110010",
      "010000" when "110011",
      "001011" when "110100",
      "000000" when "110101",
      "000000" when "110110",
      "011101" when "110111",
      "000000" when "111000",
      "000000" when "111001",
      "000000" when "111010",
      "000000" when "111011",
      "000001" when "111100",
      "000010" when "111101",
      "000000" when "111110",
      "000000" when "111111",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Subtract12_6_impl_0_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract12_6_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract12_6_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Subtract12_6_impl_0_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Subtract12_6_impl_0_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--        GenericLut_LUTData_MUX_Subtract12_6_impl_1_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract12_6_impl_1_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract12_6_impl_1_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "010101" when "000000",
      "010110" when "000001",
      "000000" when "000010",
      "000000" when "000011",
      "000000" when "000100",
      "010001" when "000101",
      "100001" when "000110",
      "010010" when "000111",
      "000000" when "001000",
      "001010" when "001001",
      "001011" when "001010",
      "000000" when "001011",
      "000000" when "001100",
      "000000" when "001101",
      "100000" when "001110",
      "001100" when "001111",
      "010011" when "010000",
      "000000" when "010001",
      "010100" when "010010",
      "011000" when "010011",
      "000000" when "010100",
      "000000" when "010101",
      "000000" when "010110",
      "000011" when "010111",
      "011001" when "011000",
      "011110" when "011001",
      "000000" when "011010",
      "000101" when "011011",
      "011111" when "011100",
      "011011" when "011101",
      "000000" when "011110",
      "000000" when "011111",
      "000000" when "100000",
      "000100" when "100001",
      "010111" when "100010",
      "000000" when "100011",
      "011010" when "100100",
      "011101" when "100101",
      "010000" when "100110",
      "000000" when "100111",
      "000000" when "101000",
      "000000" when "101001",
      "001000" when "101010",
      "001111" when "101011",
      "000000" when "101100",
      "000110" when "101101",
      "000111" when "101110",
      "001101" when "101111",
      "000000" when "110000",
      "000000" when "110001",
      "000000" when "110010",
      "001110" when "110011",
      "001001" when "110100",
      "000000" when "110101",
      "000000" when "110110",
      "011100" when "110111",
      "000000" when "111000",
      "000000" when "111001",
      "000000" when "111010",
      "000000" when "111011",
      "000001" when "111100",
      "000010" when "111101",
      "000000" when "111110",
      "000000" when "111111",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Subtract12_6_impl_1_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract12_6_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract12_6_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Subtract12_6_impl_1_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Subtract12_6_impl_1_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      Y <= s3;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      Y <= s2;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 5 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      Y <= s4;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 8 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      Y <= s7;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 7 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      Y <= s6;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      Y <= s5;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 9 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      Y <= s8;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 10 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      Y <= s9;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 26 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      Y <= s25;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 12 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      Y <= s11;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 15 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      Y <= s14;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 13 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      Y <= s12;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 30 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      Y <= s29;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      Y <= s10;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_38_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 38 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_38_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_38_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      Y <= s37;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 16 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      Y <= s15;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 31 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      Y <= s30;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 27 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      Y <= s26;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 22 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      Y <= s21;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 28 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      Y <= s27;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 21 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      Y <= s20;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 24 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      Y <= s23;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 20 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      Y <= s19;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 18 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      Y <= s17;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 29 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      Y <= s28;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 17 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      Y <= s16;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                         implementedSystem_toplevel
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity implementedSystem_toplevel is
   port ( clk, rst : in std_logic;
          x0_re_0 : in std_logic_vector(31 downto 0);
          x0_im_0 : in std_logic_vector(31 downto 0);
          x1_re_0 : in std_logic_vector(31 downto 0);
          x1_im_0 : in std_logic_vector(31 downto 0);
          x2_re_0 : in std_logic_vector(31 downto 0);
          x2_im_0 : in std_logic_vector(31 downto 0);
          x3_re_0 : in std_logic_vector(31 downto 0);
          x3_im_0 : in std_logic_vector(31 downto 0);
          x4_re_0 : in std_logic_vector(31 downto 0);
          x4_im_0 : in std_logic_vector(31 downto 0);
          x5_re_0 : in std_logic_vector(31 downto 0);
          x5_im_0 : in std_logic_vector(31 downto 0);
          x6_re_0 : in std_logic_vector(31 downto 0);
          x6_im_0 : in std_logic_vector(31 downto 0);
          x7_re_0 : in std_logic_vector(31 downto 0);
          x7_im_0 : in std_logic_vector(31 downto 0);
          x8_re_0 : in std_logic_vector(31 downto 0);
          x8_im_0 : in std_logic_vector(31 downto 0);
          x9_re_0 : in std_logic_vector(31 downto 0);
          x9_im_0 : in std_logic_vector(31 downto 0);
          x10_re_0 : in std_logic_vector(31 downto 0);
          x10_im_0 : in std_logic_vector(31 downto 0);
          x11_re_0 : in std_logic_vector(31 downto 0);
          x11_im_0 : in std_logic_vector(31 downto 0);
          x12_re_0 : in std_logic_vector(31 downto 0);
          x12_im_0 : in std_logic_vector(31 downto 0);
          x13_re_0 : in std_logic_vector(31 downto 0);
          x13_im_0 : in std_logic_vector(31 downto 0);
          x14_re_0 : in std_logic_vector(31 downto 0);
          x14_im_0 : in std_logic_vector(31 downto 0);
          x15_re_0 : in std_logic_vector(31 downto 0);
          x15_im_0 : in std_logic_vector(31 downto 0);
          y0_re_0 : out std_logic_vector(31 downto 0);
          y0_im_0 : out std_logic_vector(31 downto 0);
          y1_re_0 : out std_logic_vector(31 downto 0);
          y1_im_0 : out std_logic_vector(31 downto 0);
          y2_re_0 : out std_logic_vector(31 downto 0);
          y2_im_0 : out std_logic_vector(31 downto 0);
          y3_re_0 : out std_logic_vector(31 downto 0);
          y3_im_0 : out std_logic_vector(31 downto 0);
          y4_re_0 : out std_logic_vector(31 downto 0);
          y4_im_0 : out std_logic_vector(31 downto 0);
          y5_re_0 : out std_logic_vector(31 downto 0);
          y5_im_0 : out std_logic_vector(31 downto 0);
          y6_re_0 : out std_logic_vector(31 downto 0);
          y6_im_0 : out std_logic_vector(31 downto 0);
          y7_re_0 : out std_logic_vector(31 downto 0);
          y7_im_0 : out std_logic_vector(31 downto 0);
          y8_re_0 : out std_logic_vector(31 downto 0);
          y8_im_0 : out std_logic_vector(31 downto 0);
          y9_re_0 : out std_logic_vector(31 downto 0);
          y9_im_0 : out std_logic_vector(31 downto 0);
          y10_re_0 : out std_logic_vector(31 downto 0);
          y10_im_0 : out std_logic_vector(31 downto 0);
          y11_re_0 : out std_logic_vector(31 downto 0);
          y11_im_0 : out std_logic_vector(31 downto 0);
          y12_re_0 : out std_logic_vector(31 downto 0);
          y12_im_0 : out std_logic_vector(31 downto 0);
          y13_re_0 : out std_logic_vector(31 downto 0);
          y13_im_0 : out std_logic_vector(31 downto 0);
          y14_re_0 : out std_logic_vector(31 downto 0);
          y14_im_0 : out std_logic_vector(31 downto 0);
          y15_re_0 : out std_logic_vector(31 downto 0);
          y15_im_0 : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of implementedSystem_toplevel is
   component ModuloCounter_64_component is
      port ( clk, rst : in std_logic;
             Counter_out : out std_logic_vector(5 downto 0)   );
   end component;

   component InputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(31 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component OutputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(31 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_7_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(2 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_64_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iS_13 : in std_logic_vector(33 downto 0);
             iS_14 : in std_logic_vector(33 downto 0);
             iS_15 : in std_logic_vector(33 downto 0);
             iS_16 : in std_logic_vector(33 downto 0);
             iS_17 : in std_logic_vector(33 downto 0);
             iS_18 : in std_logic_vector(33 downto 0);
             iS_19 : in std_logic_vector(33 downto 0);
             iS_20 : in std_logic_vector(33 downto 0);
             iS_21 : in std_logic_vector(33 downto 0);
             iS_22 : in std_logic_vector(33 downto 0);
             iS_23 : in std_logic_vector(33 downto 0);
             iS_24 : in std_logic_vector(33 downto 0);
             iS_25 : in std_logic_vector(33 downto 0);
             iS_26 : in std_logic_vector(33 downto 0);
             iS_27 : in std_logic_vector(33 downto 0);
             iS_28 : in std_logic_vector(33 downto 0);
             iS_29 : in std_logic_vector(33 downto 0);
             iS_30 : in std_logic_vector(33 downto 0);
             iS_31 : in std_logic_vector(33 downto 0);
             iS_32 : in std_logic_vector(33 downto 0);
             iS_33 : in std_logic_vector(33 downto 0);
             iS_34 : in std_logic_vector(33 downto 0);
             iS_35 : in std_logic_vector(33 downto 0);
             iS_36 : in std_logic_vector(33 downto 0);
             iS_37 : in std_logic_vector(33 downto 0);
             iS_38 : in std_logic_vector(33 downto 0);
             iS_39 : in std_logic_vector(33 downto 0);
             iS_40 : in std_logic_vector(33 downto 0);
             iS_41 : in std_logic_vector(33 downto 0);
             iS_42 : in std_logic_vector(33 downto 0);
             iS_43 : in std_logic_vector(33 downto 0);
             iS_44 : in std_logic_vector(33 downto 0);
             iS_45 : in std_logic_vector(33 downto 0);
             iS_46 : in std_logic_vector(33 downto 0);
             iS_47 : in std_logic_vector(33 downto 0);
             iS_48 : in std_logic_vector(33 downto 0);
             iS_49 : in std_logic_vector(33 downto 0);
             iS_50 : in std_logic_vector(33 downto 0);
             iS_51 : in std_logic_vector(33 downto 0);
             iS_52 : in std_logic_vector(33 downto 0);
             iS_53 : in std_logic_vector(33 downto 0);
             iS_54 : in std_logic_vector(33 downto 0);
             iS_55 : in std_logic_vector(33 downto 0);
             iS_56 : in std_logic_vector(33 downto 0);
             iS_57 : in std_logic_vector(33 downto 0);
             iS_58 : in std_logic_vector(33 downto 0);
             iS_59 : in std_logic_vector(33 downto 0);
             iS_60 : in std_logic_vector(33 downto 0);
             iS_61 : in std_logic_vector(33 downto 0);
             iS_62 : in std_logic_vector(33 downto 0);
             iS_63 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(5 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_63_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iS_13 : in std_logic_vector(33 downto 0);
             iS_14 : in std_logic_vector(33 downto 0);
             iS_15 : in std_logic_vector(33 downto 0);
             iS_16 : in std_logic_vector(33 downto 0);
             iS_17 : in std_logic_vector(33 downto 0);
             iS_18 : in std_logic_vector(33 downto 0);
             iS_19 : in std_logic_vector(33 downto 0);
             iS_20 : in std_logic_vector(33 downto 0);
             iS_21 : in std_logic_vector(33 downto 0);
             iS_22 : in std_logic_vector(33 downto 0);
             iS_23 : in std_logic_vector(33 downto 0);
             iS_24 : in std_logic_vector(33 downto 0);
             iS_25 : in std_logic_vector(33 downto 0);
             iS_26 : in std_logic_vector(33 downto 0);
             iS_27 : in std_logic_vector(33 downto 0);
             iS_28 : in std_logic_vector(33 downto 0);
             iS_29 : in std_logic_vector(33 downto 0);
             iS_30 : in std_logic_vector(33 downto 0);
             iS_31 : in std_logic_vector(33 downto 0);
             iS_32 : in std_logic_vector(33 downto 0);
             iS_33 : in std_logic_vector(33 downto 0);
             iS_34 : in std_logic_vector(33 downto 0);
             iS_35 : in std_logic_vector(33 downto 0);
             iS_36 : in std_logic_vector(33 downto 0);
             iS_37 : in std_logic_vector(33 downto 0);
             iS_38 : in std_logic_vector(33 downto 0);
             iS_39 : in std_logic_vector(33 downto 0);
             iS_40 : in std_logic_vector(33 downto 0);
             iS_41 : in std_logic_vector(33 downto 0);
             iS_42 : in std_logic_vector(33 downto 0);
             iS_43 : in std_logic_vector(33 downto 0);
             iS_44 : in std_logic_vector(33 downto 0);
             iS_45 : in std_logic_vector(33 downto 0);
             iS_46 : in std_logic_vector(33 downto 0);
             iS_47 : in std_logic_vector(33 downto 0);
             iS_48 : in std_logic_vector(33 downto 0);
             iS_49 : in std_logic_vector(33 downto 0);
             iS_50 : in std_logic_vector(33 downto 0);
             iS_51 : in std_logic_vector(33 downto 0);
             iS_52 : in std_logic_vector(33 downto 0);
             iS_53 : in std_logic_vector(33 downto 0);
             iS_54 : in std_logic_vector(33 downto 0);
             iS_55 : in std_logic_vector(33 downto 0);
             iS_56 : in std_logic_vector(33 downto 0);
             iS_57 : in std_logic_vector(33 downto 0);
             iS_58 : in std_logic_vector(33 downto 0);
             iS_59 : in std_logic_vector(33 downto 0);
             iS_60 : in std_logic_vector(33 downto 0);
             iS_61 : in std_logic_vector(33 downto 0);
             iS_62 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(5 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_48_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iS_13 : in std_logic_vector(33 downto 0);
             iS_14 : in std_logic_vector(33 downto 0);
             iS_15 : in std_logic_vector(33 downto 0);
             iS_16 : in std_logic_vector(33 downto 0);
             iS_17 : in std_logic_vector(33 downto 0);
             iS_18 : in std_logic_vector(33 downto 0);
             iS_19 : in std_logic_vector(33 downto 0);
             iS_20 : in std_logic_vector(33 downto 0);
             iS_21 : in std_logic_vector(33 downto 0);
             iS_22 : in std_logic_vector(33 downto 0);
             iS_23 : in std_logic_vector(33 downto 0);
             iS_24 : in std_logic_vector(33 downto 0);
             iS_25 : in std_logic_vector(33 downto 0);
             iS_26 : in std_logic_vector(33 downto 0);
             iS_27 : in std_logic_vector(33 downto 0);
             iS_28 : in std_logic_vector(33 downto 0);
             iS_29 : in std_logic_vector(33 downto 0);
             iS_30 : in std_logic_vector(33 downto 0);
             iS_31 : in std_logic_vector(33 downto 0);
             iS_32 : in std_logic_vector(33 downto 0);
             iS_33 : in std_logic_vector(33 downto 0);
             iS_34 : in std_logic_vector(33 downto 0);
             iS_35 : in std_logic_vector(33 downto 0);
             iS_36 : in std_logic_vector(33 downto 0);
             iS_37 : in std_logic_vector(33 downto 0);
             iS_38 : in std_logic_vector(33 downto 0);
             iS_39 : in std_logic_vector(33 downto 0);
             iS_40 : in std_logic_vector(33 downto 0);
             iS_41 : in std_logic_vector(33 downto 0);
             iS_42 : in std_logic_vector(33 downto 0);
             iS_43 : in std_logic_vector(33 downto 0);
             iS_44 : in std_logic_vector(33 downto 0);
             iS_45 : in std_logic_vector(33 downto 0);
             iS_46 : in std_logic_vector(33 downto 0);
             iS_47 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(5 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_33_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iS_13 : in std_logic_vector(33 downto 0);
             iS_14 : in std_logic_vector(33 downto 0);
             iS_15 : in std_logic_vector(33 downto 0);
             iS_16 : in std_logic_vector(33 downto 0);
             iS_17 : in std_logic_vector(33 downto 0);
             iS_18 : in std_logic_vector(33 downto 0);
             iS_19 : in std_logic_vector(33 downto 0);
             iS_20 : in std_logic_vector(33 downto 0);
             iS_21 : in std_logic_vector(33 downto 0);
             iS_22 : in std_logic_vector(33 downto 0);
             iS_23 : in std_logic_vector(33 downto 0);
             iS_24 : in std_logic_vector(33 downto 0);
             iS_25 : in std_logic_vector(33 downto 0);
             iS_26 : in std_logic_vector(33 downto 0);
             iS_27 : in std_logic_vector(33 downto 0);
             iS_28 : in std_logic_vector(33 downto 0);
             iS_29 : in std_logic_vector(33 downto 0);
             iS_30 : in std_logic_vector(33 downto 0);
             iS_31 : in std_logic_vector(33 downto 0);
             iS_32 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(5 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_47_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iS_13 : in std_logic_vector(33 downto 0);
             iS_14 : in std_logic_vector(33 downto 0);
             iS_15 : in std_logic_vector(33 downto 0);
             iS_16 : in std_logic_vector(33 downto 0);
             iS_17 : in std_logic_vector(33 downto 0);
             iS_18 : in std_logic_vector(33 downto 0);
             iS_19 : in std_logic_vector(33 downto 0);
             iS_20 : in std_logic_vector(33 downto 0);
             iS_21 : in std_logic_vector(33 downto 0);
             iS_22 : in std_logic_vector(33 downto 0);
             iS_23 : in std_logic_vector(33 downto 0);
             iS_24 : in std_logic_vector(33 downto 0);
             iS_25 : in std_logic_vector(33 downto 0);
             iS_26 : in std_logic_vector(33 downto 0);
             iS_27 : in std_logic_vector(33 downto 0);
             iS_28 : in std_logic_vector(33 downto 0);
             iS_29 : in std_logic_vector(33 downto 0);
             iS_30 : in std_logic_vector(33 downto 0);
             iS_31 : in std_logic_vector(33 downto 0);
             iS_32 : in std_logic_vector(33 downto 0);
             iS_33 : in std_logic_vector(33 downto 0);
             iS_34 : in std_logic_vector(33 downto 0);
             iS_35 : in std_logic_vector(33 downto 0);
             iS_36 : in std_logic_vector(33 downto 0);
             iS_37 : in std_logic_vector(33 downto 0);
             iS_38 : in std_logic_vector(33 downto 0);
             iS_39 : in std_logic_vector(33 downto 0);
             iS_40 : in std_logic_vector(33 downto 0);
             iS_41 : in std_logic_vector(33 downto 0);
             iS_42 : in std_logic_vector(33 downto 0);
             iS_43 : in std_logic_vector(33 downto 0);
             iS_44 : in std_logic_vector(33 downto 0);
             iS_45 : in std_logic_vector(33 downto 0);
             iS_46 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(5 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_34_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iS_13 : in std_logic_vector(33 downto 0);
             iS_14 : in std_logic_vector(33 downto 0);
             iS_15 : in std_logic_vector(33 downto 0);
             iS_16 : in std_logic_vector(33 downto 0);
             iS_17 : in std_logic_vector(33 downto 0);
             iS_18 : in std_logic_vector(33 downto 0);
             iS_19 : in std_logic_vector(33 downto 0);
             iS_20 : in std_logic_vector(33 downto 0);
             iS_21 : in std_logic_vector(33 downto 0);
             iS_22 : in std_logic_vector(33 downto 0);
             iS_23 : in std_logic_vector(33 downto 0);
             iS_24 : in std_logic_vector(33 downto 0);
             iS_25 : in std_logic_vector(33 downto 0);
             iS_26 : in std_logic_vector(33 downto 0);
             iS_27 : in std_logic_vector(33 downto 0);
             iS_28 : in std_logic_vector(33 downto 0);
             iS_29 : in std_logic_vector(33 downto 0);
             iS_30 : in std_logic_vector(33 downto 0);
             iS_31 : in std_logic_vector(33 downto 0);
             iS_32 : in std_logic_vector(33 downto 0);
             iS_33 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(5 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Constant_float_8_23_1_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_0_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosnpi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinnpi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn3_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn3_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosnpi_div_2_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinnpi_div_2_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn5_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn5_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn3_mult_pi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn3_mult_pi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn7_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn7_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosnpi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinnpi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add2_5_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add2_5_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add2_6_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add2_6_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add11_6_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add11_6_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Subtract2_6_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Subtract2_6_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Subtract3_6_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Subtract3_6_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Subtract12_6_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Subtract12_6_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_38_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

signal ModCount641_out : std_logic_vector(5 downto 0) := (others => '0');
signal x0_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x0_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x1_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x1_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x2_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x2_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x3_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x3_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x4_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x4_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x5_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x5_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x6_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x6_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x7_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x7_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x8_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x8_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x9_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x9_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x10_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x10_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x11_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x11_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x12_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x12_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x13_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x13_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x14_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x14_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x15_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x15_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y0_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y0_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y1_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y1_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y2_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y2_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y3_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y3_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y4_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y4_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y5_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y5_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y6_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y6_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y7_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No14_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y7_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No15_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y8_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No16_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y8_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No17_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y9_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No18_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y9_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No19_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y10_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No20_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y10_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No21_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y11_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No22_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y11_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No23_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y12_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No24_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y12_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No25_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y13_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No26_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y13_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No27_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y14_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No28_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y14_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No29_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y15_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No30_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y15_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No31_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No32_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No33_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No34_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No35_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No36_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No37_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No38_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No39_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No40_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No41_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No42_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No43_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No44_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No45_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No46_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No47_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No48_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No49_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No50_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No51_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No52_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No53_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No54_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No55_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No56_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No57_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No58_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No59_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No60_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No61_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No62_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No63_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No64_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No65_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No66_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No67_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No68_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No69_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No70_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No71_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product31_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No72_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No73_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product31_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No74_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No75_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product31_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No76_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No77_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product31_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No78_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No79_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product31_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No80_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No81_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product31_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No82_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No83_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product31_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No84_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No85_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No86_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No87_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No88_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No89_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No90_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No91_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No92_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No93_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No94_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No95_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No96_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No97_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No98_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No99_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No100_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No101_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No102_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No103_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No104_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No105_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No106_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No107_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No108_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No109_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No110_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No111_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No112_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No113_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract3_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No114_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No115_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract3_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No116_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No117_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract6_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract6_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No118_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract6_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No119_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract6_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract6_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No120_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract6_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No121_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract10_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract10_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No122_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract10_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No123_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract12_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No124_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No125_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant2_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant11_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant4_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant13_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant5_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant14_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant6_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant15_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant7_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant16_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant8_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant17_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant9_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant18_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant1_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay76No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay76No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay76No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay76No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay76No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay76No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay77No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay77No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay77No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay77No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay77No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay77No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay77No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay44No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay44No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay44No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay44No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay44No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay44No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay44No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y0_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y0_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y1_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y1_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y2_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y2_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y3_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y3_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y4_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y4_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y5_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y5_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y6_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y6_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y7_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y7_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y8_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y8_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y9_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y9_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y10_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y10_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y11_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y11_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y12_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y12_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y13_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y13_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y14_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y14_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y15_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y15_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Add2_5_impl_0_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Add2_5_impl_1_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Add2_6_impl_0_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Add2_6_impl_1_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Add11_6_impl_0_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Add11_6_impl_1_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Subtract2_6_impl_0_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Subtract2_6_impl_1_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Subtract3_6_impl_0_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Subtract3_6_impl_1_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Subtract12_6_impl_0_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Subtract12_6_impl_1_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal SharedReg_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg360_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg408_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg434_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg463_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg465_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg470_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg477_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg481_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg483_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg485_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg500_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg508_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg510_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg512_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg528_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg531_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg533_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg534_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg536_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg582_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg587_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg588_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg592_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg601_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg602_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg604_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg605_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg607_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg616_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg620_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg626_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg629_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg634_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg644_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg646_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg649_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg666_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg667_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg670_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg676_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg680_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg681_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg682_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg688_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg690_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg702_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg703_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg705_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg706_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg721_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg724_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg725_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg731_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg736_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg740_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg745_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg750_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg751_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg756_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg757_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg761_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg762_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg763_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg765_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg771_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg774_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg775_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg823_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg844_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg864_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg869_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg870_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg873_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg874_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg875_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg877_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg878_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg879_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg880_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg881_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg890_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg891_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg892_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg893_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg894_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg895_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg896_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg897_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg898_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg905_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg915_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg919_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg923_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg925_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg930_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg944_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg945_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg946_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg949_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg950_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg951_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg952_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg953_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg954_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg955_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg956_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg958_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg959_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg960_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg961_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg962_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg963_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg964_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg965_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg966_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg967_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg969_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg970_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg971_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg972_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg973_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg974_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg975_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg976_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg977_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg978_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg979_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg980_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg981_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg982_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg983_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg984_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg985_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg986_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg987_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg988_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg989_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg990_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg991_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg992_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg993_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg994_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg995_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg996_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg997_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg999_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1000_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1001_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1002_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1003_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1004_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1005_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1006_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1007_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1008_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1009_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1010_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1012_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1013_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1014_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1015_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1016_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1017_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1018_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1019_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1020_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1021_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1022_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1023_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1024_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1025_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1026_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1028_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1029_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1030_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1031_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1032_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1033_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1034_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1035_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1036_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1038_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1039_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1040_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1041_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1042_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1043_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1044_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1045_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1046_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1047_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1048_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1049_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1050_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1051_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1052_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1053_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1054_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1055_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1056_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1058_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1059_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1060_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1061_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1062_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1064_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1065_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1066_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1067_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1068_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1069_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1070_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1071_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1072_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1073_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1074_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1075_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1077_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1078_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1079_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1080_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1081_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1082_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1083_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1084_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1085_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1087_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1088_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1089_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1090_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1091_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1092_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1093_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1094_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1095_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1096_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1097_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1098_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1099_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1100_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1101_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1102_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1105_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1127_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1128_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1130_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1132_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1133_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1138_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1142_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1143_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1144_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1145_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1146_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1147_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1148_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1149_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1150_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1151_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1153_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1154_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1155_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1156_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1157_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1159_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1160_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1161_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1162_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1163_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1164_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1165_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1166_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1167_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1168_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1169_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1170_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1171_out : std_logic_vector(33 downto 0) := (others => '0');
signal x0_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x0_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x1_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x1_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x2_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x2_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x3_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x3_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x4_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x4_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x5_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x5_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x6_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x6_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x7_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x7_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x8_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x8_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x9_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x9_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x10_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x10_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x11_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x11_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x12_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x12_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x13_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x13_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x14_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x14_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x15_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x15_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y0_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y0_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y1_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y1_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y2_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y2_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y3_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y3_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y4_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y4_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y5_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y5_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y6_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y6_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y7_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y7_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y8_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y8_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y9_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg983_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y9_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y10_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg983_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y10_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y11_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg983_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y11_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y12_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y12_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y13_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg983_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y13_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y14_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y14_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg983_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y15_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y15_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No32_out_to_Add2_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No33_out_to_Add2_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg582_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg959_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg961_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg961_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg961_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg981_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg592_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg982_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg961_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg588_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg587_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg961_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg958_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg736_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No34_out_to_Add2_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No35_out_to_Add2_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg963_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg602_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg973_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg974_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg602_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg477_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg958_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg616_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg930_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg477_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg955_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg751_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No36_out_to_Add2_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No37_out_to_Add2_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg771_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg765_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg620_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg954_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg765_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg765_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg765_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg408_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg956_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg880_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No38_out_to_Add2_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No39_out_to_Add2_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg649_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No3_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg879_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg510_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg881_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No40_out_to_Add2_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No41_out_to_Add2_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg534_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg874_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No5_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg703_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg536_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg690_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg702_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg536_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No42_out_to_Add2_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No43_out_to_Add2_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg721_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg993_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg823_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg536_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg823_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg994_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No44_out_to_Add2_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No45_out_to_Add2_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg891_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg894_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg898_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg987_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg987_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg987_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg984_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg905_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1002_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1000_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg987_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No46_out_to_Add11_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No47_out_to_Add11_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg731_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg740_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg470_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg736_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg963_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg463_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg959_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg731_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg731_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg980_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No48_out_to_Add11_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No49_out_to_Add11_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg477_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg602_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg485_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No1_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg751_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg756_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg975_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg605_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg751_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No50_out_to_Add11_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No51_out_to_Add11_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg644_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg644_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg771_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No2_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg774_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg923_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg765_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg649_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg644_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg954_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg510_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg765_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg765_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg765_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No52_out_to_Add11_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No53_out_to_Add11_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg646_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg508_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg949_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg533_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No4_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg873_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg879_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg512_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg676_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg706_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No54_out_to_Add11_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No55_out_to_Add11_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg997_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg688_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg985_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg994_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg667_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg996_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg705_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1001_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg823_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg702_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg528_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg434_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No56_out_to_Add11_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No57_out_to_Add11_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg844_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No6_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg844_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg983_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No58_out_to_Product4_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No59_out_to_Product4_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1044_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1045_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1055_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1056_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg977_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1003_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1154_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1007_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1008_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg962_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1010_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1150_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1151_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1016_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1068_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1161_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1155_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1048_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1049_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1099_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1051_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1052_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1019_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1020_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1021_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1022_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1023_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1024_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1025_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1028_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1029_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1030_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1031_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1080_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1032_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1033_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1034_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1035_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1085_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1054_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1038_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1039_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1040_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1041_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1130_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1042_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1043_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg978_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg980_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1168_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1160_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg963_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1153_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg969_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg970_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg971_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg958_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg958_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg964_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1092_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No60_out_to_Product4_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No61_out_to_Product4_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1054_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1038_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1039_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1040_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1041_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1130_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1042_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1043_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1044_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1045_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1055_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1056_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg925_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1003_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1154_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1007_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1008_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1010_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1150_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg964_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1151_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1016_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1068_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1161_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1155_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1048_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1049_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1099_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1051_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1052_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1019_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1020_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1021_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1022_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1023_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1024_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1025_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1028_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1029_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1030_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1031_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1080_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1032_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1033_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1034_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1035_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1085_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg960_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1092_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1168_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1160_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg601_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1153_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg605_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg972_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No62_out_to_Product4_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No63_out_to_Product4_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1030_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1031_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1080_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1032_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1033_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1034_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1035_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1085_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1054_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1038_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1039_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1040_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1041_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1130_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1042_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1043_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1044_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1045_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1055_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1056_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg951_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1003_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1154_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg620_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1007_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1008_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1010_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1150_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1151_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1016_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1068_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1161_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1155_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1048_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1049_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1099_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1051_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1052_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1019_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1020_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1021_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1022_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1023_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1024_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1025_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1028_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1029_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg607_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1092_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg952_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg954_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1168_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1160_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1153_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No64_out_to_Product4_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No65_out_to_Product4_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1023_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1024_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1025_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1028_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1029_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1030_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1031_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1080_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1032_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1033_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1034_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1035_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1085_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1054_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1038_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1039_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1040_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1041_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1130_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1042_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1043_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1044_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1045_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1055_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1056_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1003_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1154_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1007_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1008_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1010_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1150_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1151_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1016_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1068_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1161_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1155_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1048_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1049_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1099_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1051_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1052_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1019_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1020_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1021_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1022_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1092_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg877_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg879_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1168_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1160_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg646_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1153_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No66_out_to_Product4_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No67_out_to_Product4_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1048_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1049_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1099_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1051_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1052_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1019_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1020_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1021_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1022_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1023_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1024_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1025_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1028_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1029_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1030_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1031_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1080_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1032_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1033_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1034_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1035_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1085_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1054_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1038_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1039_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1040_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1041_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1130_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1042_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1043_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1044_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1045_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1055_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1056_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1003_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1154_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1007_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1008_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1010_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1150_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1151_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1016_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1068_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1161_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1155_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg945_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1092_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg680_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg682_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1168_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1160_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg667_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg667_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1153_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No68_out_to_Product4_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No69_out_to_Product4_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg892_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1151_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1016_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1068_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1161_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1155_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1048_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1049_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1099_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1051_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1052_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1019_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1020_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1021_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1022_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1023_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1024_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1025_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1028_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1029_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1030_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1031_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1080_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1032_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1033_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1034_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1035_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1085_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1054_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1038_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1039_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1040_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1041_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1130_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1042_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1043_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1044_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1045_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1055_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1056_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1003_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1154_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg688_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1007_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1008_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg690_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1010_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1150_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1153_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg893_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg870_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg688_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1092_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg724_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1168_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1160_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No70_out_to_Product4_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No71_out_to_Product4_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1154_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg688_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1007_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1008_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1010_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1150_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg994_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1151_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1016_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1068_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1161_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1155_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1048_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1049_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1099_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1051_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1052_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1019_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1020_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1021_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1022_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1023_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1024_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1025_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1028_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1029_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1030_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1031_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1080_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1032_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1033_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1034_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1035_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1085_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1054_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1038_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1039_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1040_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1041_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1130_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1042_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1043_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1044_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1045_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1055_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1056_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg999_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1003_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1160_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg989_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg890_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg892_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1153_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg995_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg894_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg895_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg984_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg990_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg896_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1092_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1000_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1168_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No72_out_to_Product31_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No73_out_to_Product31_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1094_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1105_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1046_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1170_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1004_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1166_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1006_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1171_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1060_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1013_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1014_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1015_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1017_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1018_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1047_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1049_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1050_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1051_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1156_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1072_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg958_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1074_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg958_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1077_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1029_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1159_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1081_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1082_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1084_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1036_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1089_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1090_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1145_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1091_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1132_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1133_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1093_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg980_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg958_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1061_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1062_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg963_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1067_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1097_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg971_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg971_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1101_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1070_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1071_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1073_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1075_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg965_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1079_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1083_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1087_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1088_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No74_out_to_Product31_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No75_out_to_Product31_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1089_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1090_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1145_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1091_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1132_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1133_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1094_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1105_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1046_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1170_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1004_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1166_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1006_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1171_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1060_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg601_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1013_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1014_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1015_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1017_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1018_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1047_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1049_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1050_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1051_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1156_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1072_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1074_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1077_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1029_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1159_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1081_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1082_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1084_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1036_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1087_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1088_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg960_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1093_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1061_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1062_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg965_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1067_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1097_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg604_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg919_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg919_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1101_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1070_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1071_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1073_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1075_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg601_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1079_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1083_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg972_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No76_out_to_Product31_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No77_out_to_Product31_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1159_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1081_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1082_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1084_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1036_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1089_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1090_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1145_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1091_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1132_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1133_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1094_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1105_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1046_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1170_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1004_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1166_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1006_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1171_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1060_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1013_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1014_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1015_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1017_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1018_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1047_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1049_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1050_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1051_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1156_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1072_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1074_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1077_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1029_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1079_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1083_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg607_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1087_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1088_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1093_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg954_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1061_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1062_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1067_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1097_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg629_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg944_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg944_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1101_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1070_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1071_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1073_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1075_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No78_out_to_Product31_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No79_out_to_Product31_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1074_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1077_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1029_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1159_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1081_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1082_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1084_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1036_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1089_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1090_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1145_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1091_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1132_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1133_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1094_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1105_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1046_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1170_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1004_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1166_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1006_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1171_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1060_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1013_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1014_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1015_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1017_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1018_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1047_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1049_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1050_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1051_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1156_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1072_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1073_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1075_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1079_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1083_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1087_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1088_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1093_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg879_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg644_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1061_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1062_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg646_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg646_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1067_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1097_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg869_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1101_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1070_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1071_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No80_out_to_Product31_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No81_out_to_Product31_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1049_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1050_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1051_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1156_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1072_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1074_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1077_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1029_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1159_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1081_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1082_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1084_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1036_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1089_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1090_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1145_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1091_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1132_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1133_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1094_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1105_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1046_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1170_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1004_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1166_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1006_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1171_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1060_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1013_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1014_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1015_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1017_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1018_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1047_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1097_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1101_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1070_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1071_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1073_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1075_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1079_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1083_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg945_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1087_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1088_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1093_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg682_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1061_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1062_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg646_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg667_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg667_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1067_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No82_out_to_Product31_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No83_out_to_Product31_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1013_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1014_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1015_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1017_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1018_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1047_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1049_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1050_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1051_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1156_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1072_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1074_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1077_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1029_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1159_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1081_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1082_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1084_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1036_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1089_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1090_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1145_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1091_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1132_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1133_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1094_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1105_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1046_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1170_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1004_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1166_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1006_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1171_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1060_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1067_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1097_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1101_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1070_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1071_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1073_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1075_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1079_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1083_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg870_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1087_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1088_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg688_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1093_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1061_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1062_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg667_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No84_out_to_Product31_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No85_out_to_Product31_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1166_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1006_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1171_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1060_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg890_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1013_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1014_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1015_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1017_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1018_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1047_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1049_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1050_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1051_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1156_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1072_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg984_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1074_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1077_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1029_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1159_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1081_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1082_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1084_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1036_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1089_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1090_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1145_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1091_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1132_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1133_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1094_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1105_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1046_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1170_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1004_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1061_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1062_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg989_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1067_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1097_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg895_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1101_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1070_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1071_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1073_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1075_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1079_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1083_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg896_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1087_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1088_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg984_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1093_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1000_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No86_out_to_Subtract2_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No87_out_to_Subtract2_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg582_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg959_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg963_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg961_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg731_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay44No_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg731_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg360_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg961_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg745_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg736_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg958_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg465_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No88_out_to_Subtract2_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No89_out_to_Subtract2_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg963_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg602_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg973_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg483_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg761_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg958_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg751_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg751_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay44No1_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg750_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No1_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg763_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No90_out_to_Subtract2_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No91_out_to_Subtract2_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg620_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg771_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg765_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg765_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg765_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg954_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg500_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay44No2_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg775_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No2_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No92_out_to_Subtract2_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No93_out_to_Subtract2_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg510_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg649_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg531_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg649_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg508_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg953_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg879_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg508_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No10_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay44No3_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg510_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay77No3_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No4_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No94_out_to_Subtract2_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No95_out_to_Subtract2_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg873_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg873_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg703_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No5_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg690_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg878_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg702_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay44No4_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No12_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay76No4_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No96_out_to_Subtract2_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No97_out_to_Subtract2_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg997_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg985_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg667_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg996_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay77No5_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg536_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg823_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay44No5_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No98_out_to_Subtract2_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No99_out_to_Subtract2_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg993_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg434_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg994_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg994_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg706_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1001_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg823_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No100_out_to_Product32_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No101_out_to_Product32_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1149_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1055_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1056_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1170_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1005_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1059_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg961_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1009_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1169_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1167_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1012_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1065_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1014_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1016_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1068_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1069_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1097_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1098_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg971_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1100_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg966_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1053_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1102_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1162_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1157_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1026_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg965_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1078_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1165_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1127_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg962_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1128_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1054_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1144_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1130_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1146_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1148_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg979_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg976_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1095_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1058_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1171_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1060_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg965_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg960_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg961_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1064_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1066_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1096_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1099_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg971_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1101_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg967_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg958_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1163_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg958_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1164_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1077_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg964_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1079_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1138_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg965_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg966_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg961_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1142_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1143_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg958_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg958_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg959_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg962_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1147_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No102_out_to_Product32_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No103_out_to_Product32_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1054_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1144_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1130_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1146_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1149_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1055_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1056_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1170_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1005_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1059_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1009_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1169_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1167_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1012_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1065_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1014_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1016_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1068_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1069_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1097_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1098_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg919_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1100_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg915_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1053_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1102_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1162_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1157_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1026_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg601_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1078_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1165_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1127_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1128_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1142_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1143_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1147_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1148_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1095_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1058_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1171_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1060_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1064_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg605_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1066_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1096_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg604_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1099_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg919_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1101_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg958_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1163_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1164_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1077_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1079_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1138_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg915_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No104_out_to_Product32_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No105_out_to_Product32_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1165_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1127_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1128_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1054_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1144_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1130_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1146_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1149_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1055_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1056_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1170_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1005_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1059_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1009_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1169_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1167_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1012_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1065_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1014_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1016_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1068_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1069_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1097_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1098_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg944_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1100_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1053_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1102_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1162_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1157_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1026_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1078_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1079_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1138_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg626_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1142_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1143_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1147_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1148_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg953_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg950_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1095_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1058_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1171_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1060_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1064_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1066_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1096_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg629_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1099_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg944_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1101_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1163_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg620_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1164_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1077_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No106_out_to_Product32_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No107_out_to_Product32_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1157_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1026_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1078_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1165_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1127_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1128_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1054_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1144_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1130_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1146_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1149_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1055_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1056_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1170_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1005_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1059_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1009_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1169_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1167_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1012_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1065_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1014_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1016_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1068_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1069_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1097_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1098_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg869_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1100_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg864_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1053_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1102_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1162_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1163_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1164_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1077_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1079_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1138_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg644_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1142_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1143_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1147_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1148_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg878_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg875_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1095_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1058_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1171_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1060_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg644_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1064_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1066_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1096_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1099_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1101_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No108_out_to_Product32_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No109_out_to_Product32_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1097_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1098_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1100_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg670_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1053_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1102_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1162_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1157_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1026_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1078_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1165_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1127_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg666_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1128_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1054_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1144_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1130_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1146_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1149_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1055_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1056_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1170_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1005_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1059_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1009_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1169_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1167_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1012_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1065_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1014_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1016_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1068_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1069_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1099_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1101_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1163_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1164_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1077_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1079_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1138_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg864_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1142_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1143_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg666_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1147_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1148_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg681_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1095_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1058_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1171_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1060_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg644_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg688_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1064_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1066_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1096_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No110_out_to_Product32_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No111_out_to_Product32_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1012_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1065_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1014_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1016_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1068_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1069_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1097_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1098_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1100_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1053_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1102_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1162_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1157_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1026_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg690_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1078_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1165_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1127_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1128_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1054_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1144_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1130_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1146_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1149_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1055_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1056_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1170_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1005_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1059_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1009_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1169_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1167_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1066_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1096_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1099_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1101_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1163_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg688_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1164_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1077_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1079_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1138_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg670_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg690_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1142_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1143_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1147_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1148_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg725_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1095_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1058_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1171_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1060_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg890_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1064_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No112_out_to_Product32_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No113_out_to_Product32_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1005_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1059_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1009_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1169_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1167_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1012_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1065_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1014_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1016_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1068_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1069_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1097_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1098_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg895_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1100_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg992_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1053_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1102_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1162_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1157_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1026_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1078_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1165_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1127_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg988_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1128_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1054_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg983_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg983_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1144_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1130_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1146_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1149_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1055_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1056_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg983_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1170_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1171_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1060_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg991_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1064_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg894_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg892_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1066_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1096_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1099_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1101_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg993_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1163_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg983_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg984_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1164_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1077_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg990_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1079_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1138_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg991_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg992_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg987_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1142_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1143_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg984_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg988_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg984_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1147_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1148_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1095_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1058_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No114_out_to_Subtract3_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No115_out_to_Subtract3_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg646_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg644_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg676_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No11_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay76No3_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay77No4_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No116_out_to_Subtract3_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No117_out_to_Subtract3_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg721_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg897_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg989_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg987_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg984_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No6_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay44No6_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg844_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1000_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg984_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No118_out_to_Subtract6_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No119_out_to_Subtract6_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg477_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg602_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg974_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg974_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg602_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg605_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg477_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg634_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg774_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg750_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg762_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No8_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg757_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay76No1_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay77No1_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg955_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No120_out_to_Subtract6_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No121_out_to_Subtract6_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg644_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg946_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg765_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg765_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg771_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg771_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No9_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg765_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay76No2_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay77No2_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg771_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg880_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No3_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No122_out_to_Subtract10_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No123_out_to_Subtract10_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg960_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg963_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No7_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg958_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg981_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay76No_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay77No_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg588_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg588_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg980_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg958_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_60_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg756_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_61_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_62_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg750_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_63_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg481_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_64_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No124_out_to_Subtract12_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No125_out_to_Subtract12_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg891_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg894_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg986_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay43No13_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay76No6_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay77No6_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg983_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   ModCount641_instance: ModuloCounter_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Counter_out => ModCount641_out);
x0_re_0_IEEE <= x0_re_0;
   x0_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x0_re_0_out,
                 X => x0_re_0_IEEE);
x0_im_0_IEEE <= x0_im_0;
   x0_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x0_im_0_out,
                 X => x0_im_0_IEEE);
x1_re_0_IEEE <= x1_re_0;
   x1_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x1_re_0_out,
                 X => x1_re_0_IEEE);
x1_im_0_IEEE <= x1_im_0;
   x1_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x1_im_0_out,
                 X => x1_im_0_IEEE);
x2_re_0_IEEE <= x2_re_0;
   x2_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x2_re_0_out,
                 X => x2_re_0_IEEE);
x2_im_0_IEEE <= x2_im_0;
   x2_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x2_im_0_out,
                 X => x2_im_0_IEEE);
x3_re_0_IEEE <= x3_re_0;
   x3_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x3_re_0_out,
                 X => x3_re_0_IEEE);
x3_im_0_IEEE <= x3_im_0;
   x3_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x3_im_0_out,
                 X => x3_im_0_IEEE);
x4_re_0_IEEE <= x4_re_0;
   x4_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x4_re_0_out,
                 X => x4_re_0_IEEE);
x4_im_0_IEEE <= x4_im_0;
   x4_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x4_im_0_out,
                 X => x4_im_0_IEEE);
x5_re_0_IEEE <= x5_re_0;
   x5_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x5_re_0_out,
                 X => x5_re_0_IEEE);
x5_im_0_IEEE <= x5_im_0;
   x5_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x5_im_0_out,
                 X => x5_im_0_IEEE);
x6_re_0_IEEE <= x6_re_0;
   x6_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x6_re_0_out,
                 X => x6_re_0_IEEE);
x6_im_0_IEEE <= x6_im_0;
   x6_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x6_im_0_out,
                 X => x6_im_0_IEEE);
x7_re_0_IEEE <= x7_re_0;
   x7_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x7_re_0_out,
                 X => x7_re_0_IEEE);
x7_im_0_IEEE <= x7_im_0;
   x7_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x7_im_0_out,
                 X => x7_im_0_IEEE);
x8_re_0_IEEE <= x8_re_0;
   x8_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x8_re_0_out,
                 X => x8_re_0_IEEE);
x8_im_0_IEEE <= x8_im_0;
   x8_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x8_im_0_out,
                 X => x8_im_0_IEEE);
x9_re_0_IEEE <= x9_re_0;
   x9_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x9_re_0_out,
                 X => x9_re_0_IEEE);
x9_im_0_IEEE <= x9_im_0;
   x9_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x9_im_0_out,
                 X => x9_im_0_IEEE);
x10_re_0_IEEE <= x10_re_0;
   x10_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x10_re_0_out,
                 X => x10_re_0_IEEE);
x10_im_0_IEEE <= x10_im_0;
   x10_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x10_im_0_out,
                 X => x10_im_0_IEEE);
x11_re_0_IEEE <= x11_re_0;
   x11_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x11_re_0_out,
                 X => x11_re_0_IEEE);
x11_im_0_IEEE <= x11_im_0;
   x11_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x11_im_0_out,
                 X => x11_im_0_IEEE);
x12_re_0_IEEE <= x12_re_0;
   x12_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x12_re_0_out,
                 X => x12_re_0_IEEE);
x12_im_0_IEEE <= x12_im_0;
   x12_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x12_im_0_out,
                 X => x12_im_0_IEEE);
x13_re_0_IEEE <= x13_re_0;
   x13_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x13_re_0_out,
                 X => x13_re_0_IEEE);
x13_im_0_IEEE <= x13_im_0;
   x13_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x13_im_0_out,
                 X => x13_im_0_IEEE);
x14_re_0_IEEE <= x14_re_0;
   x14_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x14_re_0_out,
                 X => x14_re_0_IEEE);
x14_im_0_IEEE <= x14_im_0;
   x14_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x14_im_0_out,
                 X => x14_im_0_IEEE);
x15_re_0_IEEE <= x15_re_0;
   x15_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x15_re_0_out,
                 X => x15_re_0_IEEE);
x15_im_0_IEEE <= x15_im_0;
   x15_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x15_im_0_out,
                 X => x15_im_0_IEEE);
   y0_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y0_re_0_IEEE,
                 X => Delay1No_out);
y0_re_0 <= y0_re_0_IEEE;

SharedReg36_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg36_out;
SharedReg62_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg62_out;
SharedReg234_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg234_out;
SharedReg260_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg260_out;
SharedReg114_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg114_out;
SharedReg139_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg139_out;
SharedReg310_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg310_out;
   MUX_y0_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg36_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg62_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg234_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg260_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg114_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg139_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg310_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y0_re_0_0_LUT_out,
                 oMux => MUX_y0_re_0_0_out);

   Delay1No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y0_re_0_0_out,
                 Y => Delay1No_out);
   y0_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y0_im_0_IEEE,
                 X => Delay1No1_out);
y0_im_0 <= y0_im_0_IEEE;

SharedReg208_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg208_out;
SharedReg234_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg234_out;
SharedReg88_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg88_out;
SharedReg114_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg114_out;
SharedReg285_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg285_out;
SharedReg310_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg310_out;
SharedReg163_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg163_out;
   MUX_y0_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg208_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg234_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg88_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg114_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg285_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg310_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg163_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y0_im_0_0_LUT_out,
                 oMux => MUX_y0_im_0_0_out);

   Delay1No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y0_im_0_0_out,
                 Y => Delay1No1_out);
   y1_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y1_re_0_IEEE,
                 X => Delay1No2_out);
y1_re_0 <= y1_re_0_IEEE;

SharedReg36_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg36_out;
SharedReg62_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg62_out;
SharedReg234_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg234_out;
SharedReg260_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg260_out;
SharedReg285_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg285_out;
SharedReg310_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg310_out;
SharedReg186_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg186_out;
   MUX_y1_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg36_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg62_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg234_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg260_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg285_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg310_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg186_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y1_re_0_0_LUT_out,
                 oMux => MUX_y1_re_0_0_out);

   Delay1No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y1_re_0_0_out,
                 Y => Delay1No2_out);
   y1_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y1_im_0_IEEE,
                 X => Delay1No3_out);
y1_im_0 <= y1_im_0_IEEE;

SharedReg208_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg208_out;
SharedReg234_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg234_out;
SharedReg88_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg88_out;
SharedReg114_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg114_out;
SharedReg139_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg139_out;
SharedReg163_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg163_out;
SharedReg332_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg332_out;
   MUX_y1_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg208_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg234_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg88_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg114_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg139_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg163_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg332_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y1_im_0_0_LUT_out,
                 oMux => MUX_y1_im_0_0_out);

   Delay1No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y1_im_0_0_out,
                 Y => Delay1No3_out);
   y2_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y2_re_0_IEEE,
                 X => Delay1No4_out);
y2_re_0 <= y2_re_0_IEEE;

SharedReg36_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg36_out;
SharedReg62_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg62_out;
SharedReg88_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg88_out;
SharedReg114_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg114_out;
SharedReg285_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg285_out;
SharedReg310_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg310_out;
SharedReg186_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg186_out;
   MUX_y2_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg36_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg62_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg88_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg114_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg285_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg310_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg186_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y2_re_0_0_LUT_out,
                 oMux => MUX_y2_re_0_0_out);

   Delay1No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y2_re_0_0_out,
                 Y => Delay1No4_out);
   y2_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y2_im_0_IEEE,
                 X => Delay1No5_out);
y2_im_0 <= y2_im_0_IEEE;

SharedReg208_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg208_out;
SharedReg234_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg234_out;
SharedReg260_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg260_out;
SharedReg285_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg285_out;
SharedReg139_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg139_out;
SharedReg163_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg163_out;
SharedReg332_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg332_out;
   MUX_y2_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg208_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg234_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg260_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg285_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg139_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg163_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg332_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y2_im_0_0_LUT_out,
                 oMux => MUX_y2_im_0_0_out);

   Delay1No5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y2_im_0_0_out,
                 Y => Delay1No5_out);
   y3_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y3_re_0_IEEE,
                 X => Delay1No6_out);
y3_re_0 <= y3_re_0_IEEE;

SharedReg36_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg36_out;
SharedReg208_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg208_out;
SharedReg234_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg234_out;
SharedReg260_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg260_out;
SharedReg285_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg285_out;
SharedReg310_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg310_out;
SharedReg186_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg186_out;
   MUX_y3_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg36_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg208_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg234_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg260_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg285_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg310_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg186_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y3_re_0_0_LUT_out,
                 oMux => MUX_y3_re_0_0_out);

   Delay1No6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y3_re_0_0_out,
                 Y => Delay1No6_out);
   y3_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y3_im_0_IEEE,
                 X => Delay1No7_out);
y3_im_0 <= y3_im_0_IEEE;

SharedReg36_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg36_out;
SharedReg208_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg208_out;
SharedReg234_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg234_out;
SharedReg260_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg260_out;
SharedReg285_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg285_out;
SharedReg310_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg310_out;
SharedReg163_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg163_out;
   MUX_y3_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg36_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg208_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg234_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg260_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg285_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg310_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg163_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y3_im_0_0_LUT_out,
                 oMux => MUX_y3_im_0_0_out);

   Delay1No7_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y3_im_0_0_out,
                 Y => Delay1No7_out);
   y4_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y4_re_0_IEEE,
                 X => Delay1No8_out);
y4_re_0 <= y4_re_0_IEEE;

SharedReg36_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg36_out;
SharedReg62_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg62_out;
SharedReg62_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg62_out;
SharedReg88_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg88_out;
SharedReg260_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg260_out;
SharedReg285_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg285_out;
SharedReg310_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg310_out;
   MUX_y4_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg36_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg62_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg62_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg88_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg260_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg285_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg310_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y4_re_0_0_LUT_out,
                 oMux => MUX_y4_re_0_0_out);

   Delay1No8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y4_re_0_0_out,
                 Y => Delay1No8_out);
   y4_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y4_im_0_IEEE,
                 X => Delay1No9_out);
y4_im_0 <= y4_im_0_IEEE;

SharedReg208_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg208_out;
SharedReg234_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg234_out;
SharedReg234_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg234_out;
SharedReg260_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg260_out;
SharedReg114_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg114_out;
SharedReg139_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg139_out;
SharedReg163_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg163_out;
   MUX_y4_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg208_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg234_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg234_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg260_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg114_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg139_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg163_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y4_im_0_0_LUT_out,
                 oMux => MUX_y4_im_0_0_out);

   Delay1No9_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y4_im_0_0_out,
                 Y => Delay1No9_out);
   y5_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y5_re_0_IEEE,
                 X => Delay1No10_out);
y5_re_0 <= y5_re_0_IEEE;

SharedReg36_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg36_out;
SharedReg62_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg62_out;
SharedReg234_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg234_out;
SharedReg260_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg260_out;
SharedReg285_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg285_out;
SharedReg310_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg310_out;
SharedReg163_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg163_out;
   MUX_y5_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg36_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg62_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg234_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg260_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg285_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg310_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg163_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y5_re_0_0_LUT_out,
                 oMux => MUX_y5_re_0_0_out);

   Delay1No10_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y5_re_0_0_out,
                 Y => Delay1No10_out);
   y5_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y5_im_0_IEEE,
                 X => Delay1No11_out);
y5_im_0 <= y5_im_0_IEEE;

SharedReg36_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg36_out;
SharedReg208_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg208_out;
SharedReg62_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg62_out;
SharedReg88_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg88_out;
SharedReg114_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg114_out;
SharedReg139_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg139_out;
SharedReg163_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg163_out;
   MUX_y5_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg36_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg208_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg62_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg88_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg114_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg139_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg163_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y5_im_0_0_LUT_out,
                 oMux => MUX_y5_im_0_0_out);

   Delay1No11_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y5_im_0_0_out,
                 Y => Delay1No11_out);
   y6_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y6_re_0_IEEE,
                 X => Delay1No12_out);
y6_re_0 <= y6_re_0_IEEE;

SharedReg36_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg36_out;
SharedReg62_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg62_out;
SharedReg88_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg88_out;
SharedReg114_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg114_out;
SharedReg285_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg285_out;
SharedReg310_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg310_out;
SharedReg186_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg186_out;
   MUX_y6_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg36_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg62_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg88_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg114_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg285_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg310_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg186_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y6_re_0_0_LUT_out,
                 oMux => MUX_y6_re_0_0_out);

   Delay1No12_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y6_re_0_0_out,
                 Y => Delay1No12_out);
   y6_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y6_im_0_IEEE,
                 X => Delay1No13_out);
y6_im_0 <= y6_im_0_IEEE;

SharedReg36_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg36_out;
SharedReg62_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg62_out;
SharedReg88_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg88_out;
SharedReg114_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg114_out;
SharedReg285_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg285_out;
SharedReg310_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg310_out;
SharedReg163_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg163_out;
   MUX_y6_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg36_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg62_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg88_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg114_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg285_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg310_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg163_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y6_im_0_0_LUT_out,
                 oMux => MUX_y6_im_0_0_out);

   Delay1No13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y6_im_0_0_out,
                 Y => Delay1No13_out);
   y7_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y7_re_0_IEEE,
                 X => Delay1No14_out);
y7_re_0 <= y7_re_0_IEEE;

SharedReg208_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg208_out;
SharedReg62_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg62_out;
SharedReg88_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg88_out;
SharedReg114_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg114_out;
SharedReg139_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg139_out;
SharedReg163_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg163_out;
SharedReg186_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg186_out;
   MUX_y7_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg208_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg62_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg88_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg114_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg139_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg163_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg186_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y7_re_0_0_LUT_out,
                 oMux => MUX_y7_re_0_0_out);

   Delay1No14_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y7_re_0_0_out,
                 Y => Delay1No14_out);
   y7_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y7_im_0_IEEE,
                 X => Delay1No15_out);
y7_im_0 <= y7_im_0_IEEE;

SharedReg36_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg36_out;
SharedReg208_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg208_out;
SharedReg234_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg234_out;
SharedReg260_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg260_out;
SharedReg285_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg285_out;
SharedReg310_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg310_out;
SharedReg310_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg310_out;
   MUX_y7_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg36_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg208_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg234_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg260_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg285_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg310_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg310_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y7_im_0_0_LUT_out,
                 oMux => MUX_y7_im_0_0_out);

   Delay1No15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y7_im_0_0_out,
                 Y => Delay1No15_out);
   y8_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y8_re_0_IEEE,
                 X => Delay1No16_out);
y8_re_0 <= y8_re_0_IEEE;

SharedReg567_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg567_out;
SharedReg593_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg593_out;
SharedReg906_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg906_out;
SharedReg931_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg931_out;
SharedReg640_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg640_out;
SharedReg661_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg661_out;
SharedReg685_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg685_out;
   MUX_y8_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg567_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg593_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg906_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg931_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg640_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg661_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg685_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y8_re_0_0_LUT_out,
                 oMux => MUX_y8_re_0_0_out);

   Delay1No16_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y8_re_0_0_out,
                 Y => Delay1No16_out);
   y8_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y8_im_0_IEEE,
                 X => Delay1No17_out);
y8_im_0 <= y8_im_0_IEEE;

SharedReg957_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg957_out;
SharedReg906_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg906_out;
SharedReg617_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg617_out;
SharedReg640_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg640_out;
SharedReg855_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg855_out;
SharedReg685_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg685_out;
SharedReg707_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg707_out;
   MUX_y8_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg957_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg906_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg617_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg640_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg855_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg685_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg707_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y8_im_0_0_LUT_out,
                 oMux => MUX_y8_im_0_0_out);

   Delay1No17_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y8_im_0_0_out,
                 Y => Delay1No17_out);
   y9_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y9_re_0_IEEE,
                 X => Delay1No18_out);
y9_re_0 <= y9_re_0_IEEE;

SharedReg957_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg957_out;
SharedReg906_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg906_out;
SharedReg617_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg617_out;
SharedReg640_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg640_out;
SharedReg661_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg661_out;
SharedReg707_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg707_out;
SharedReg983_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg983_out;
   MUX_y9_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg957_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg906_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg617_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg640_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg661_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg707_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg983_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y9_re_0_0_LUT_out,
                 oMux => MUX_y9_re_0_0_out);

   Delay1No18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y9_re_0_0_out,
                 Y => Delay1No18_out);
   y9_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y9_im_0_IEEE,
                 X => Delay1No19_out);
y9_im_0 <= y9_im_0_IEEE;

SharedReg957_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg957_out;
SharedReg906_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg906_out;
SharedReg617_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg617_out;
SharedReg640_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg640_out;
SharedReg661_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg661_out;
SharedReg707_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg707_out;
SharedReg707_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg707_out;
   MUX_y9_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg957_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg906_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg617_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg640_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg661_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg707_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg707_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y9_im_0_0_LUT_out,
                 oMux => MUX_y9_im_0_0_out);

   Delay1No19_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y9_im_0_0_out,
                 Y => Delay1No19_out);
   y10_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y10_re_0_IEEE,
                 X => Delay1No20_out);
y10_re_0 <= y10_re_0_IEEE;

SharedReg957_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg957_out;
SharedReg906_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg906_out;
SharedReg931_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg931_out;
SharedReg855_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg855_out;
SharedReg661_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg661_out;
SharedReg707_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg707_out;
SharedReg983_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg983_out;
   MUX_y10_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg957_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg906_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg931_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg855_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg661_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg707_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg983_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y10_re_0_0_LUT_out,
                 oMux => MUX_y10_re_0_0_out);

   Delay1No20_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y10_re_0_0_out,
                 Y => Delay1No20_out);
   y10_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y10_im_0_IEEE,
                 X => Delay1No21_out);
y10_im_0 <= y10_im_0_IEEE;

SharedReg567_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg567_out;
SharedReg593_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg593_out;
SharedReg617_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg617_out;
SharedReg640_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg640_out;
SharedReg855_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg855_out;
SharedReg685_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg685_out;
SharedReg882_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg882_out;
   MUX_y10_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg567_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg593_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg617_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg640_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg855_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg685_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg882_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y10_im_0_0_LUT_out,
                 oMux => MUX_y10_im_0_0_out);

   Delay1No21_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y10_im_0_0_out,
                 Y => Delay1No21_out);
   y11_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y11_re_0_IEEE,
                 X => Delay1No22_out);
y11_re_0 <= y11_re_0_IEEE;

SharedReg957_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg957_out;
SharedReg593_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg593_out;
SharedReg617_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg617_out;
SharedReg640_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg640_out;
SharedReg661_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg661_out;
SharedReg707_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg707_out;
SharedReg983_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg983_out;
   MUX_y11_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg957_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg593_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg617_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg640_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg661_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg707_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg983_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y11_re_0_0_LUT_out,
                 oMux => MUX_y11_re_0_0_out);

   Delay1No22_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y11_re_0_0_out,
                 Y => Delay1No22_out);
   y11_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y11_im_0_IEEE,
                 X => Delay1No23_out);
y11_im_0 <= y11_im_0_IEEE;

SharedReg567_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg567_out;
SharedReg957_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg957_out;
SharedReg906_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg906_out;
SharedReg931_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg931_out;
SharedReg855_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg855_out;
SharedReg685_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg685_out;
SharedReg707_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg707_out;
   MUX_y11_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg567_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg957_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg906_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg931_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg855_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg685_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg707_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y11_im_0_0_LUT_out,
                 oMux => MUX_y11_im_0_0_out);

   Delay1No23_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y11_im_0_0_out,
                 Y => Delay1No23_out);
   y12_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y12_re_0_IEEE,
                 X => Delay1No24_out);
y12_re_0 <= y12_re_0_IEEE;

SharedReg957_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg957_out;
SharedReg906_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg906_out;
SharedReg906_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg906_out;
SharedReg931_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg931_out;
SharedReg640_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg640_out;
SharedReg661_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg661_out;
SharedReg707_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg707_out;
   MUX_y12_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg957_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg906_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg906_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg931_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg640_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg661_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg707_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y12_re_0_0_LUT_out,
                 oMux => MUX_y12_re_0_0_out);

   Delay1No24_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y12_re_0_0_out,
                 Y => Delay1No24_out);
   y12_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y12_im_0_IEEE,
                 X => Delay1No25_out);
y12_im_0 <= y12_im_0_IEEE;

SharedReg567_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg567_out;
SharedReg593_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg593_out;
SharedReg593_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg593_out;
SharedReg617_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg617_out;
SharedReg931_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg931_out;
SharedReg855_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg855_out;
SharedReg685_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg685_out;
   MUX_y12_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg567_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg593_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg593_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg617_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg931_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg855_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg685_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y12_im_0_0_LUT_out,
                 oMux => MUX_y12_im_0_0_out);

   Delay1No25_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y12_im_0_0_out,
                 Y => Delay1No25_out);
   y13_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y13_re_0_IEEE,
                 X => Delay1No26_out);
y13_re_0 <= y13_re_0_IEEE;

SharedReg957_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg957_out;
SharedReg593_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg593_out;
SharedReg906_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg906_out;
SharedReg931_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg931_out;
SharedReg640_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg640_out;
SharedReg661_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg661_out;
SharedReg983_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg983_out;
   MUX_y13_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg957_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg593_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg906_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg931_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg640_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg661_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg983_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y13_re_0_0_LUT_out,
                 oMux => MUX_y13_re_0_0_out);

   Delay1No26_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y13_re_0_0_out,
                 Y => Delay1No26_out);
   y13_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y13_im_0_IEEE,
                 X => Delay1No27_out);
y13_im_0 <= y13_im_0_IEEE;

SharedReg567_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg567_out;
SharedReg957_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg957_out;
SharedReg906_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg906_out;
SharedReg931_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg931_out;
SharedReg855_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg855_out;
SharedReg685_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg685_out;
SharedReg882_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg882_out;
   MUX_y13_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg567_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg957_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg906_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg931_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg855_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg685_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg882_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y13_im_0_0_LUT_out,
                 oMux => MUX_y13_im_0_0_out);

   Delay1No27_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y13_im_0_0_out,
                 Y => Delay1No27_out);
   y14_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y14_re_0_IEEE,
                 X => Delay1No28_out);
y14_re_0 <= y14_re_0_IEEE;

SharedReg567_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg567_out;
SharedReg593_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg593_out;
SharedReg617_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg617_out;
SharedReg931_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg931_out;
SharedReg640_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg640_out;
SharedReg661_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg661_out;
SharedReg882_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg882_out;
   MUX_y14_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg567_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg593_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg617_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg931_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg640_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg661_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg882_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y14_re_0_0_LUT_out,
                 oMux => MUX_y14_re_0_0_out);

   Delay1No28_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y14_re_0_0_out,
                 Y => Delay1No28_out);
   y14_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y14_im_0_IEEE,
                 X => Delay1No29_out);
y14_im_0 <= y14_im_0_IEEE;

SharedReg983_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg983_out;
SharedReg957_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg957_out;
SharedReg906_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg906_out;
SharedReg931_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg931_out;
SharedReg640_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg640_out;
SharedReg855_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg855_out;
SharedReg685_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg685_out;
   MUX_y14_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg983_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg957_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg906_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg931_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg640_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg855_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg685_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y14_im_0_0_LUT_out,
                 oMux => MUX_y14_im_0_0_out);

   Delay1No29_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y14_im_0_0_out,
                 Y => Delay1No29_out);
   y15_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y15_re_0_IEEE,
                 X => Delay1No30_out);
y15_re_0 <= y15_re_0_IEEE;

SharedReg957_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg957_out;
SharedReg593_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg593_out;
SharedReg617_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg617_out;
SharedReg640_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg640_out;
SharedReg661_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg661_out;
SharedReg707_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg707_out;
SharedReg882_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg882_out;
   MUX_y15_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg957_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg593_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg617_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg640_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg661_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg707_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg882_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y15_re_0_0_LUT_out,
                 oMux => MUX_y15_re_0_0_out);

   Delay1No30_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y15_re_0_0_out,
                 Y => Delay1No30_out);
   y15_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y15_im_0_IEEE,
                 X => Delay1No31_out);
y15_im_0 <= y15_im_0_IEEE;

SharedReg957_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg957_out;
SharedReg593_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg593_out;
SharedReg617_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg617_out;
SharedReg640_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg640_out;
SharedReg661_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg661_out;
SharedReg707_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg707_out;
SharedReg707_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg707_out;
   MUX_y15_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg957_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg593_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg617_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg640_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg661_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg707_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg707_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y15_im_0_0_LUT_out,
                 oMux => MUX_y15_im_0_0_out);

   Delay1No31_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y15_im_0_0_out,
                 Y => Delay1No31_out);

Delay1No32_out_to_Add2_0_impl_parent_implementedSystem_port_0_cast <= Delay1No32_out;
Delay1No33_out_to_Add2_0_impl_parent_implementedSystem_port_1_cast <= Delay1No33_out;
   Add2_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_0_impl_out,
                 X => Delay1No32_out_to_Add2_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No33_out_to_Add2_0_impl_parent_implementedSystem_port_1_cast);

SharedReg41_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg41_out;
SharedReg_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg_out;
SharedReg2_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg2_out;
SharedReg5_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg5_out;
SharedReg4_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg7_out;
SharedReg10_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg10_out;
SharedReg9_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg9_out;
SharedReg13_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg13_out;
SharedReg356_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg356_out;
SharedReg356_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg356_out;
SharedReg45_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg45_out;
SharedReg582_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg582_out;
SharedReg466_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg466_out;
SharedReg457_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg457_out;
SharedReg746_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg746_out;
SharedReg350_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg350_out;
SharedReg350_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg350_out;
SharedReg55_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg55_out;
SharedReg356_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg356_out;
SharedReg585_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg585_out;
SharedReg959_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg959_out;
SharedReg569_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg569_out;
SharedReg229_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg229_out;
SharedReg570_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg570_out;
SharedReg961_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg961_out;
SharedReg212_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg212_out;
SharedReg350_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg350_out;
SharedReg213_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_29_cast <= SharedReg213_out;
SharedReg358_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_30_cast <= SharedReg358_out;
SharedReg567_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_31_cast <= SharedReg567_out;
SharedReg968_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_32_cast <= SharedReg968_out;
SharedReg961_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_33_cast <= SharedReg961_out;
SharedReg208_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_34_cast <= SharedReg208_out;
SharedReg576_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_35_cast <= SharedReg576_out;
SharedReg569_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_36_cast <= SharedReg569_out;
SharedReg53_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_37_cast <= SharedReg53_out;
SharedReg364_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_38_cast <= SharedReg364_out;
SharedReg461_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_39_cast <= SharedReg461_out;
SharedReg459_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_40_cast <= SharedReg459_out;
SharedReg917_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_41_cast <= SharedReg917_out;
SharedReg350_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_42_cast <= SharedReg350_out;
SharedReg54_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_43_cast <= SharedReg54_out;
SharedReg568_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_44_cast <= SharedReg568_out;
SharedReg568_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_45_cast <= SharedReg568_out;
SharedReg38_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_46_cast <= SharedReg38_out;
SharedReg584_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_47_cast <= SharedReg584_out;
SharedReg961_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_48_cast <= SharedReg961_out;
SharedReg213_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_49_cast <= SharedReg213_out;
SharedReg41_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_50_cast <= SharedReg41_out;
SharedReg350_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_51_cast <= SharedReg350_out;
SharedReg41_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_52_cast <= SharedReg41_out;
SharedReg573_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_53_cast <= SharedReg573_out;
SharedReg573_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_54_cast <= SharedReg573_out;
SharedReg361_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_55_cast <= SharedReg361_out;
SharedReg350_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_56_cast <= SharedReg350_out;
SharedReg573_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_57_cast <= SharedReg573_out;
SharedReg215_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_58_cast <= SharedReg215_out;
SharedReg217_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_59_cast <= SharedReg217_out;
SharedReg576_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_60_cast <= SharedReg576_out;
SharedReg734_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_61_cast <= SharedReg734_out;
SharedReg364_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_62_cast <= SharedReg364_out;
SharedReg352_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_63_cast <= SharedReg352_out;
SharedReg352_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_64_cast <= SharedReg352_out;
   MUX_Add2_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg41_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg356_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg45_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg582_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg466_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg457_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg746_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg350_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg350_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg55_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg356_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg2_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg585_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg959_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg569_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg229_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg570_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg961_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg212_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg350_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg213_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg358_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg5_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg567_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg968_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg961_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg208_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg576_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg569_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg53_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg364_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg461_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg459_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg4_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg917_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg350_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg54_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg568_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg568_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg38_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg584_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg961_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg213_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg41_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg7_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg350_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg41_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg573_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg573_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg361_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg350_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg573_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg215_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg217_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg576_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg10_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg734_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg364_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg352_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg352_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg9_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg13_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg356_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add2_0_impl_0_out);

   Delay1No32_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_0_impl_0_out,
                 Y => Delay1No32_out);

SharedReg40_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg40_out;
SharedReg18_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg20_out;
SharedReg23_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg23_out;
SharedReg22_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg25_out;
SharedReg28_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg28_out;
SharedReg27_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg27_out;
SharedReg31_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg31_out;
SharedReg462_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg462_out;
SharedReg459_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg459_out;
SharedReg46_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg46_out;
SharedReg581_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg581_out;
SharedReg363_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg363_out;
SharedReg729_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg729_out;
SharedReg359_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg359_out;
SharedReg455_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg455_out;
SharedReg357_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg357_out;
SharedReg36_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg36_out;
SharedReg455_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg455_out;
SharedReg569_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg569_out;
SharedReg591_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg591_out;
SharedReg981_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg981_out;
SharedReg213_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg213_out;
SharedReg592_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg592_out;
SharedReg982_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg982_out;
SharedReg233_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg233_out;
SharedReg461_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg461_out;
SharedReg208_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_29_cast <= SharedReg208_out;
SharedReg350_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_30_cast <= SharedReg350_out;
SharedReg572_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_31_cast <= SharedReg572_out;
SharedReg567_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_32_cast <= SharedReg567_out;
SharedReg571_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_33_cast <= SharedReg571_out;
SharedReg210_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_34_cast <= SharedReg210_out;
SharedReg567_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_35_cast <= SharedReg567_out;
SharedReg961_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_36_cast <= SharedReg961_out;
SharedReg208_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_37_cast <= SharedReg208_out;
SharedReg357_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_38_cast <= SharedReg357_out;
SharedReg734_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_39_cast <= SharedReg734_out;
SharedReg733_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_40_cast <= SharedReg733_out;
SharedReg593_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_41_cast <= SharedReg593_out;
SharedReg456_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_42_cast <= SharedReg456_out;
SharedReg36_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_43_cast <= SharedReg36_out;
SharedReg588_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_44_cast <= SharedReg588_out;
SharedReg587_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_45_cast <= SharedReg587_out;
SharedReg227_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_46_cast <= SharedReg227_out;
SharedReg961_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_47_cast <= SharedReg961_out;
SharedReg590_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_48_cast <= SharedReg590_out;
SharedReg59_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_49_cast <= SharedReg59_out;
SharedReg231_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_50_cast <= SharedReg231_out;
SharedReg457_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_51_cast <= SharedReg457_out;
SharedReg208_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_52_cast <= SharedReg208_out;
SharedReg567_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_53_cast <= SharedReg567_out;
SharedReg958_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_54_cast <= SharedReg958_out;
SharedReg455_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_55_cast <= SharedReg455_out;
SharedReg457_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_56_cast <= SharedReg457_out;
SharedReg567_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_57_cast <= SharedReg567_out;
SharedReg209_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_58_cast <= SharedReg209_out;
SharedReg208_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_59_cast <= SharedReg208_out;
SharedReg568_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_60_cast <= SharedReg568_out;
SharedReg736_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_61_cast <= SharedReg736_out;
SharedReg459_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_62_cast <= SharedReg459_out;
SharedReg455_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_63_cast <= SharedReg455_out;
SharedReg455_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_64_cast <= SharedReg455_out;
   MUX_Add2_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg40_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg18_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg459_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg46_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg581_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg363_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg729_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg359_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg455_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg357_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg36_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg455_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg20_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg569_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg591_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg981_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg213_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg592_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg982_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg233_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg461_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg208_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg350_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg23_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg572_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg567_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg571_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg210_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg567_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg961_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg208_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg357_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg734_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg733_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg22_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg593_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg456_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg36_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg588_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg587_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg227_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg961_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg590_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg59_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg231_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg25_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg457_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg208_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg567_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg958_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg455_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg457_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg567_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg209_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg208_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg568_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg28_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg736_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg459_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg455_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg455_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg27_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg31_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg462_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add2_0_impl_1_out);

   Delay1No33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_0_impl_1_out,
                 Y => Delay1No33_out);

Delay1No34_out_to_Add2_1_impl_parent_implementedSystem_port_0_cast <= Delay1No34_out;
Delay1No35_out_to_Add2_1_impl_parent_implementedSystem_port_1_cast <= Delay1No35_out;
   Add2_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_1_impl_out,
                 X => Delay1No34_out_to_Add2_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No35_out_to_Add2_1_impl_parent_implementedSystem_port_1_cast);

SharedReg365_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg365_out;
SharedReg963_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg963_out;
SharedReg69_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg69_out;
SharedReg243_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg243_out;
SharedReg602_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg602_out;
SharedReg752_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg752_out;
SharedReg379_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg379_out;
SharedReg367_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg367_out;
SharedReg367_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg367_out;
SharedReg213_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg213_out;
SharedReg_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg_out;
SharedReg2_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg2_out;
SharedReg5_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg5_out;
SharedReg4_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg7_out;
SharedReg10_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg10_out;
SharedReg9_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg9_out;
SharedReg13_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg13_out;
SharedReg371_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg371_out;
SharedReg371_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg371_out;
SharedReg71_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg71_out;
SharedReg973_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg973_out;
SharedReg482_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg482_out;
SharedReg473_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg473_out;
SharedReg764_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg764_out;
SharedReg365_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg365_out;
SharedReg365_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg365_out;
SharedReg747_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg747_out;
SharedReg371_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_29_cast <= SharedReg371_out;
SharedReg974_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_30_cast <= SharedReg974_out;
SharedReg908_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_31_cast <= SharedReg908_out;
SharedReg595_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_32_cast <= SharedReg595_out;
SharedReg81_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_33_cast <= SharedReg81_out;
SharedReg596_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_34_cast <= SharedReg596_out;
SharedReg910_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_35_cast <= SharedReg910_out;
SharedReg238_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_36_cast <= SharedReg238_out;
SharedReg365_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_37_cast <= SharedReg365_out;
SharedReg67_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_38_cast <= SharedReg67_out;
SharedReg373_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_39_cast <= SharedReg373_out;
SharedReg234_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_40_cast <= SharedReg234_out;
SharedReg619_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_41_cast <= SharedReg619_out;
SharedReg246_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_42_cast <= SharedReg246_out;
SharedReg234_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_43_cast <= SharedReg234_out;
SharedReg602_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_44_cast <= SharedReg602_out;
SharedReg595_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_45_cast <= SharedReg595_out;
SharedReg78_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_46_cast <= SharedReg78_out;
SharedReg379_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_47_cast <= SharedReg379_out;
SharedReg477_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_48_cast <= SharedReg477_out;
SharedReg475_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_49_cast <= SharedReg475_out;
SharedReg942_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_50_cast <= SharedReg942_out;
SharedReg621_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_51_cast <= SharedReg621_out;
SharedReg79_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_52_cast <= SharedReg79_out;
SharedReg594_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_53_cast <= SharedReg594_out;
SharedReg594_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_54_cast <= SharedReg594_out;
SharedReg365_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_55_cast <= SharedReg365_out;
SharedReg372_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_56_cast <= SharedReg372_out;
SharedReg471_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_57_cast <= SharedReg471_out;
SharedReg597_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_58_cast <= SharedReg597_out;
SharedReg471_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_59_cast <= SharedReg471_out;
SharedReg380_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_60_cast <= SharedReg380_out;
SharedReg753_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_61_cast <= SharedReg753_out;
SharedReg239_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_62_cast <= SharedReg239_out;
SharedReg754_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_63_cast <= SharedReg754_out;
SharedReg236_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_64_cast <= SharedReg236_out;
   MUX_Add2_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg365_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg963_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg2_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg5_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg4_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg7_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg10_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg9_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg13_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg371_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg371_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg69_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg71_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg973_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg482_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg473_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg764_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg365_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg365_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg747_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg371_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg974_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg243_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg908_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg595_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg81_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg596_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg910_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg238_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg365_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg67_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg373_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg234_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg602_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg619_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg246_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg234_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg602_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg595_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg78_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg379_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg477_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg475_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg942_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg752_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg621_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg79_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg594_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg594_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg365_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg372_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg471_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg597_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg471_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg380_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg379_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg753_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg239_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg754_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg236_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg367_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg367_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg213_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add2_1_impl_0_out);

   Delay1No34_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_1_impl_0_out,
                 Y => Delay1No34_out);

SharedReg473_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg473_out;
SharedReg957_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg957_out;
SharedReg63_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg63_out;
SharedReg62_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg62_out;
SharedReg958_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg958_out;
SharedReg754_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg754_out;
SharedReg475_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg475_out;
SharedReg471_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg471_out;
SharedReg471_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg471_out;
SharedReg66_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg66_out;
SharedReg18_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg20_out;
SharedReg23_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg23_out;
SharedReg22_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg25_out;
SharedReg28_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg28_out;
SharedReg27_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg27_out;
SharedReg31_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg31_out;
SharedReg478_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg478_out;
SharedReg475_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg475_out;
SharedReg72_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg72_out;
SharedReg608_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg608_out;
SharedReg378_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg378_out;
SharedReg747_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg747_out;
SharedReg374_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg374_out;
SharedReg471_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg471_out;
SharedReg372_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg372_out;
SharedReg478_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg478_out;
SharedReg471_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_29_cast <= SharedReg471_out;
SharedReg595_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_30_cast <= SharedReg595_out;
SharedReg615_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_31_cast <= SharedReg615_out;
SharedReg929_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_32_cast <= SharedReg929_out;
SharedReg239_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_33_cast <= SharedReg239_out;
SharedReg616_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_34_cast <= SharedReg616_out;
SharedReg930_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_35_cast <= SharedReg930_out;
SharedReg259_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_36_cast <= SharedReg259_out;
SharedReg477_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_37_cast <= SharedReg477_out;
SharedReg234_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_38_cast <= SharedReg234_out;
SharedReg365_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_39_cast <= SharedReg365_out;
SharedReg240_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_40_cast <= SharedReg240_out;
SharedReg955_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_41_cast <= SharedReg955_out;
SharedReg62_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_42_cast <= SharedReg62_out;
SharedReg236_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_43_cast <= SharedReg236_out;
SharedReg593_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_44_cast <= SharedReg593_out;
SharedReg910_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_45_cast <= SharedReg910_out;
SharedReg208_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_46_cast <= SharedReg208_out;
SharedReg372_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_47_cast <= SharedReg372_out;
SharedReg752_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_48_cast <= SharedReg752_out;
SharedReg751_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_49_cast <= SharedReg751_out;
SharedReg617_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_50_cast <= SharedReg617_out;
SharedReg910_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_51_cast <= SharedReg910_out;
SharedReg62_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_52_cast <= SharedReg62_out;
SharedReg612_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_53_cast <= SharedReg612_out;
SharedReg611_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_54_cast <= SharedReg611_out;
SharedReg749_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_55_cast <= SharedReg749_out;
SharedReg365_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_56_cast <= SharedReg365_out;
SharedReg755_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_57_cast <= SharedReg755_out;
SharedReg928_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_58_cast <= SharedReg928_out;
SharedReg747_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_59_cast <= SharedReg747_out;
SharedReg488_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_60_cast <= SharedReg488_out;
SharedReg747_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_61_cast <= SharedReg747_out;
SharedReg62_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_62_cast <= SharedReg62_out;
SharedReg366_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_63_cast <= SharedReg366_out;
SharedReg106_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_64_cast <= SharedReg106_out;
   MUX_Add2_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg473_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg957_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg18_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg20_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg23_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg22_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg25_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg28_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg27_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg31_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg478_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg475_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg63_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg72_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg608_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg378_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg747_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg374_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg471_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg372_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg478_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg471_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg595_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg62_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg615_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg929_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg239_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg616_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg930_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg259_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg477_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg234_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg365_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg240_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg958_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg955_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg62_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg236_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg593_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg910_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg208_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg372_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg752_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg751_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg617_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg754_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg910_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg62_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg612_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg611_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg749_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg365_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg755_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg928_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg747_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg488_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg475_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg747_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg62_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg366_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg106_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg471_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg471_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg66_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add2_1_impl_1_out);

   Delay1No35_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_1_impl_1_out,
                 Y => Delay1No35_out);

Delay1No36_out_to_Add2_2_impl_parent_implementedSystem_port_0_cast <= Delay1No36_out;
Delay1No37_out_to_Add2_2_impl_parent_implementedSystem_port_1_cast <= Delay1No37_out;
   Add2_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_2_impl_out,
                 X => Delay1No36_out_to_Add2_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No37_out_to_Add2_2_impl_parent_implementedSystem_port_1_cast);

SharedReg387_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg387_out;
SharedReg487_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg487_out;
SharedReg910_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg910_out;
SharedReg487_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg487_out;
SharedReg395_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg395_out;
SharedReg771_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg771_out;
SharedReg92_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg92_out;
SharedReg772_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg772_out;
SharedReg262_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg262_out;
SharedReg380_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg380_out;
SharedReg599_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg599_out;
SharedReg241_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg241_out;
SharedReg96_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg96_out;
SharedReg916_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg916_out;
SharedReg770_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg770_out;
SharedReg394_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg394_out;
SharedReg382_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg382_out;
SharedReg382_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg382_out;
SharedReg239_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg239_out;
SharedReg_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg_out;
SharedReg2_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg2_out;
SharedReg5_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg5_out;
SharedReg4_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg7_out;
SharedReg10_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg10_out;
SharedReg9_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg9_out;
SharedReg13_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg13_out;
SharedReg773_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg773_out;
SharedReg386_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_29_cast <= SharedReg386_out;
SharedReg96_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_30_cast <= SharedReg96_out;
SharedReg921_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_31_cast <= SharedReg921_out;
SharedReg498_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_32_cast <= SharedReg498_out;
SharedReg489_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_33_cast <= SharedReg489_out;
SharedReg782_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_34_cast <= SharedReg782_out;
SharedReg380_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_35_cast <= SharedReg380_out;
SharedReg380_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_36_cast <= SharedReg380_out;
SharedReg765_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_37_cast <= SharedReg765_out;
SharedReg386_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_38_cast <= SharedReg386_out;
SharedReg922_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_39_cast <= SharedReg922_out;
SharedReg262_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_40_cast <= SharedReg262_out;
SharedReg514_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_41_cast <= SharedReg514_out;
SharedReg380_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_42_cast <= SharedReg380_out;
SharedReg620_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_43_cast <= SharedReg620_out;
SharedReg935_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_44_cast <= SharedReg935_out;
SharedReg264_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_45_cast <= SharedReg264_out;
SharedReg380_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_46_cast <= SharedReg380_out;
SharedReg92_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_47_cast <= SharedReg92_out;
SharedReg388_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_48_cast <= SharedReg388_out;
SharedReg260_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_49_cast <= SharedReg260_out;
SharedReg642_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_50_cast <= SharedReg642_out;
SharedReg133_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_51_cast <= SharedReg133_out;
SharedReg260_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_52_cast <= SharedReg260_out;
SharedReg627_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_53_cast <= SharedReg627_out;
SharedReg619_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_54_cast <= SharedReg619_out;
SharedReg630_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_55_cast <= SharedReg630_out;
SharedReg502_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_56_cast <= SharedReg502_out;
SharedReg386_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_57_cast <= SharedReg386_out;
SharedReg640_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_58_cast <= SharedReg640_out;
SharedReg794_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_59_cast <= SharedReg794_out;
SharedReg297_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_60_cast <= SharedReg297_out;
SharedReg380_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_61_cast <= SharedReg380_out;
SharedReg89_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_62_cast <= SharedReg89_out;
SharedReg380_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_63_cast <= SharedReg380_out;
SharedReg277_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_64_cast <= SharedReg277_out;
   MUX_Add2_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg387_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg487_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg599_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg241_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg96_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg916_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg770_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg394_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg382_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg382_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg239_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg910_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg2_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg5_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg4_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg7_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg10_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg9_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg13_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg773_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg386_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg96_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg487_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg921_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg498_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg489_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg782_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg380_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg380_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg765_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg386_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg922_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg262_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg395_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg514_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg380_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg620_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg935_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg264_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg380_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg92_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg388_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg260_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg642_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg771_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg133_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg260_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg627_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg619_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg630_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg502_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg386_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg640_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg794_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg297_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg92_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg380_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg89_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg380_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg277_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg772_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg262_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg380_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add2_2_impl_0_out);

   Delay1No36_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_2_impl_0_out,
                 Y => Delay1No36_out);

SharedReg380_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg380_out;
SharedReg773_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg773_out;
SharedReg954_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg954_out;
SharedReg765_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg765_out;
SharedReg504_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg504_out;
SharedReg765_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg765_out;
SharedReg88_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg88_out;
SharedReg381_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg381_out;
SharedReg131_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg131_out;
SharedReg489_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg489_out;
SharedReg906_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg906_out;
SharedReg89_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg89_out;
SharedReg88_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg88_out;
SharedReg907_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg907_out;
SharedReg772_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg772_out;
SharedReg491_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg491_out;
SharedReg487_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg487_out;
SharedReg487_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg487_out;
SharedReg91_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg91_out;
SharedReg18_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg20_out;
SharedReg23_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg23_out;
SharedReg22_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg25_out;
SharedReg28_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg28_out;
SharedReg27_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg27_out;
SharedReg31_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg31_out;
SharedReg495_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg495_out;
SharedReg491_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_29_cast <= SharedReg491_out;
SharedReg97_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_30_cast <= SharedReg97_out;
SharedReg632_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_31_cast <= SharedReg632_out;
SharedReg393_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_32_cast <= SharedReg393_out;
SharedReg765_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_33_cast <= SharedReg765_out;
SharedReg389_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_34_cast <= SharedReg389_out;
SharedReg487_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_35_cast <= SharedReg487_out;
SharedReg387_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_36_cast <= SharedReg387_out;
SharedReg494_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_37_cast <= SharedReg494_out;
SharedReg487_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_38_cast <= SharedReg487_out;
SharedReg619_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_39_cast <= SharedReg619_out;
SharedReg113_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_40_cast <= SharedReg113_out;
SharedReg408_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_41_cast <= SharedReg408_out;
SharedReg488_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_42_cast <= SharedReg488_out;
SharedReg639_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_43_cast <= SharedReg639_out;
SharedReg956_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_44_cast <= SharedReg956_out;
SharedReg284_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_45_cast <= SharedReg284_out;
SharedReg493_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_46_cast <= SharedReg493_out;
SharedReg88_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_47_cast <= SharedReg88_out;
SharedReg380_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_48_cast <= SharedReg380_out;
SharedReg266_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_49_cast <= SharedReg266_out;
SharedReg880_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_50_cast <= SharedReg880_out;
SharedReg265_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_51_cast <= SharedReg265_out;
SharedReg262_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_52_cast <= SharedReg262_out;
SharedReg617_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_53_cast <= SharedReg617_out;
SharedReg935_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_54_cast <= SharedReg935_out;
SharedReg593_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_55_cast <= SharedReg593_out;
SharedReg770_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_56_cast <= SharedReg770_out;
SharedReg384_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_57_cast <= SharedReg384_out;
SharedReg645_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_58_cast <= SharedReg645_out;
SharedReg784_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_59_cast <= SharedReg784_out;
SharedReg260_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_60_cast <= SharedReg260_out;
SharedReg767_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_61_cast <= SharedReg767_out;
SharedReg110_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_62_cast <= SharedReg110_out;
SharedReg488_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_63_cast <= SharedReg488_out;
SharedReg88_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_64_cast <= SharedReg88_out;
   MUX_Add2_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg380_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg773_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg906_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg89_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg88_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg907_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg772_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg491_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg487_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg487_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg91_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg18_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg954_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg20_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg23_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg22_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg25_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg28_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg27_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg31_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg495_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg491_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg97_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg765_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg632_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg393_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg765_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg389_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg487_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg387_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg494_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg487_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg619_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg113_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg504_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg408_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg488_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg639_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg956_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg284_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg493_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg88_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg380_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg266_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg880_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg765_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg265_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg262_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg617_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg935_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg593_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg770_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg384_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg645_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg784_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg260_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg88_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg767_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg110_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg488_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg88_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg381_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg131_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg489_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add2_2_impl_1_out);

   Delay1No37_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_2_impl_1_out,
                 Y => Delay1No37_out);

Delay1No38_out_to_Add2_3_impl_parent_implementedSystem_port_0_cast <= Delay1No38_out;
Delay1No39_out_to_Add2_3_impl_parent_implementedSystem_port_1_cast <= Delay1No39_out;
   Add2_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_3_impl_out,
                 X => Delay1No38_out_to_Add2_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No39_out_to_Add2_3_impl_parent_implementedSystem_port_1_cast);

SharedReg518_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg518_out;
SharedReg401_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg401_out;
SharedReg855_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg855_out;
SharedReg812_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg812_out;
SharedReg320_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg320_out;
SharedReg395_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg395_out;
SharedReg115_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg115_out;
SharedReg395_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg395_out;
SharedReg128_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg128_out;
SharedReg402_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg402_out;
SharedReg503_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg503_out;
SharedReg935_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg935_out;
SharedReg503_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg503_out;
SharedReg410_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg410_out;
SharedReg789_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg789_out;
SharedReg118_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg118_out;
SharedReg790_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg790_out;
SharedReg287_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg287_out;
SharedReg395_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg395_out;
SharedReg623_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg623_out;
SharedReg267_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg267_out;
SharedReg122_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg122_out;
SharedReg941_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg941_out;
SharedReg788_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg788_out;
SharedReg409_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg409_out;
SharedReg397_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg397_out;
SharedReg397_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg397_out;
SharedReg785_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg785_out;
SharedReg_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_29_cast <= SharedReg_out;
SharedReg2_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_30_cast <= SharedReg2_out;
SharedReg5_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_31_cast <= SharedReg5_out;
SharedReg4_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_32_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_33_cast <= SharedReg7_out;
SharedReg10_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_34_cast <= SharedReg10_out;
SharedReg9_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_35_cast <= SharedReg9_out;
SharedReg13_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_36_cast <= SharedReg13_out;
SharedReg791_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_37_cast <= SharedReg791_out;
SharedReg401_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_38_cast <= SharedReg401_out;
SharedReg122_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_39_cast <= SharedReg122_out;
SharedReg649_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_40_cast <= SharedReg649_out;
SharedReg4_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_41_cast <= SharedReg4_out;
Delay43No3_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_42_cast <= Delay43No3_out;
SharedReg800_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_43_cast <= SharedReg800_out;
SharedReg395_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_44_cast <= SharedReg395_out;
SharedReg395_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_45_cast <= SharedReg395_out;
SharedReg783_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_46_cast <= SharedReg783_out;
SharedReg401_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_47_cast <= SharedReg401_out;
SharedReg948_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_48_cast <= SharedReg948_out;
SharedReg116_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_49_cast <= SharedReg116_out;
SharedReg530_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_50_cast <= SharedReg530_out;
SharedReg521_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_51_cast <= SharedReg521_out;
SharedReg643_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_52_cast <= SharedReg643_out;
SharedReg859_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_53_cast <= SharedReg859_out;
SharedReg289_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_54_cast <= SharedReg289_out;
SharedReg304_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_55_cast <= SharedReg304_out;
SharedReg395_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_56_cast <= SharedReg395_out;
SharedReg505_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_57_cast <= SharedReg505_out;
SharedReg857_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_58_cast <= SharedReg857_out;
SharedReg141_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_59_cast <= SharedReg141_out;
SharedReg410_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_60_cast <= SharedReg410_out;
SharedReg650_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_61_cast <= SharedReg650_out;
SharedReg125_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_62_cast <= SharedReg125_out;
SharedReg125_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_63_cast <= SharedReg125_out;
SharedReg410_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_64_cast <= SharedReg410_out;
   MUX_Add2_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg518_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg401_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg503_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg935_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg503_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg410_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg789_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg118_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg790_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg287_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg395_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg623_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg855_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg267_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg122_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg941_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg788_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg409_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg397_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg397_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg785_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg2_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg812_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg5_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg4_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg7_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg10_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg9_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg13_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg791_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg401_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg122_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg649_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg320_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg4_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => Delay43No3_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg800_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg395_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg395_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg783_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg401_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg948_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg116_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg530_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg395_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg521_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg643_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg859_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg289_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg304_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg395_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg505_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg857_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg141_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg410_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg115_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg650_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg125_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg125_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg410_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg395_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg128_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg402_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add2_3_impl_0_out);

   Delay1No38_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_3_impl_0_out,
                 Y => Delay1No38_out);

SharedReg788_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg788_out;
SharedReg399_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg399_out;
SharedReg860_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg860_out;
SharedReg802_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg802_out;
SharedReg114_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg114_out;
SharedReg785_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg785_out;
SharedReg135_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg135_out;
SharedReg504_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg504_out;
SharedReg114_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg114_out;
SharedReg395_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg395_out;
SharedReg791_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg791_out;
SharedReg879_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg879_out;
SharedReg783_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg783_out;
SharedReg520_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg520_out;
SharedReg783_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg783_out;
SharedReg114_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg114_out;
SharedReg396_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg396_out;
SharedReg154_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg154_out;
SharedReg505_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg505_out;
SharedReg931_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg931_out;
SharedReg115_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg115_out;
SharedReg114_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg114_out;
SharedReg932_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg932_out;
SharedReg790_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg790_out;
SharedReg507_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg507_out;
SharedReg503_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg503_out;
SharedReg503_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg503_out;
SharedReg784_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg784_out;
SharedReg18_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_29_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_30_cast <= SharedReg20_out;
SharedReg23_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_31_cast <= SharedReg23_out;
SharedReg22_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_32_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_33_cast <= SharedReg25_out;
SharedReg28_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_34_cast <= SharedReg28_out;
SharedReg27_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_35_cast <= SharedReg27_out;
SharedReg31_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_36_cast <= SharedReg31_out;
SharedReg511_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_37_cast <= SharedReg511_out;
SharedReg507_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_38_cast <= SharedReg507_out;
SharedReg123_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_39_cast <= SharedReg123_out;
SharedReg650_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_40_cast <= SharedReg650_out;
SharedReg22_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_41_cast <= SharedReg22_out;
SharedReg514_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_42_cast <= SharedReg514_out;
SharedReg404_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_43_cast <= SharedReg404_out;
SharedReg503_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_44_cast <= SharedReg503_out;
SharedReg402_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_45_cast <= SharedReg402_out;
SharedReg510_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_46_cast <= SharedReg510_out;
SharedReg503_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_47_cast <= SharedReg503_out;
SharedReg619_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_48_cast <= SharedReg619_out;
SharedReg138_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_49_cast <= SharedReg138_out;
SharedReg423_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_50_cast <= SharedReg423_out;
SharedReg801_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_51_cast <= SharedReg801_out;
SharedReg660_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_52_cast <= SharedReg660_out;
SharedReg881_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_53_cast <= SharedReg881_out;
SharedReg309_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_54_cast <= SharedReg309_out;
SharedReg114_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_55_cast <= SharedReg114_out;
SharedReg787_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_56_cast <= SharedReg787_out;
SharedReg783_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_57_cast <= SharedReg783_out;
SharedReg683_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_58_cast <= SharedReg683_out;
SharedReg330_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_59_cast <= SharedReg330_out;
SharedReg520_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_60_cast <= SharedReg520_out;
SharedReg640_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_61_cast <= SharedReg640_out;
SharedReg114_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_62_cast <= SharedReg114_out;
SharedReg261_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_63_cast <= SharedReg261_out;
SharedReg525_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_64_cast <= SharedReg525_out;
   MUX_Add2_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg788_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg399_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg791_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg879_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg783_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg520_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg783_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg114_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg396_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg154_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg505_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg931_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg860_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg115_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg114_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg932_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg790_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg507_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg503_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg503_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg784_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg18_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg20_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg802_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg23_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg22_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg25_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg28_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg27_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg31_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg511_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg507_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg123_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg650_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg114_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg22_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg514_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg404_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg503_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg402_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg510_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg503_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg619_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg138_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg423_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg785_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg801_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg660_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg881_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg309_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg114_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg787_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg783_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg683_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg330_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg520_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg135_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg640_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg114_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg261_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg525_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg504_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg114_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg395_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add2_3_impl_1_out);

   Delay1No39_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_3_impl_1_out,
                 Y => Delay1No39_out);

Delay1No40_out_to_Add2_4_impl_parent_implementedSystem_port_0_cast <= Delay1No40_out;
Delay1No41_out_to_Add2_4_impl_parent_implementedSystem_port_1_cast <= Delay1No41_out;
   Add2_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_4_impl_out,
                 X => Delay1No40_out_to_Add2_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No41_out_to_Add2_4_impl_parent_implementedSystem_port_1_cast);

SharedReg410_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg410_out;
SharedReg521_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg521_out;
SharedReg663_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg663_out;
SharedReg312_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg312_out;
SharedReg425_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg425_out;
SharedReg672_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg672_out;
SharedReg150_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg150_out;
SharedReg150_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg150_out;
SharedReg425_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg425_out;
SharedReg534_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg534_out;
SharedReg416_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg416_out;
SharedReg685_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg685_out;
SharedReg830_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg830_out;
SharedReg174_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg174_out;
SharedReg410_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg410_out;
SharedReg140_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg140_out;
SharedReg410_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg410_out;
SharedReg302_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg302_out;
SharedReg417_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg417_out;
SharedReg519_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg519_out;
SharedReg859_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg859_out;
SharedReg519_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg519_out;
SharedReg425_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg425_out;
SharedReg807_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg807_out;
SharedReg142_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg142_out;
SharedReg808_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg808_out;
SharedReg312_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg312_out;
SharedReg872_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg872_out;
SharedReg937_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_29_cast <= SharedReg937_out;
SharedReg292_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_30_cast <= SharedReg292_out;
SharedReg146_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_31_cast <= SharedReg146_out;
SharedReg865_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_32_cast <= SharedReg865_out;
SharedReg806_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_33_cast <= SharedReg806_out;
SharedReg424_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_34_cast <= SharedReg424_out;
SharedReg412_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_35_cast <= SharedReg412_out;
SharedReg412_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_36_cast <= SharedReg412_out;
SharedReg803_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_37_cast <= SharedReg803_out;
SharedReg_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_38_cast <= SharedReg_out;
SharedReg2_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_39_cast <= SharedReg2_out;
SharedReg17_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_40_cast <= SharedReg17_out;
SharedReg695_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_41_cast <= SharedReg695_out;
SharedReg11_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_42_cast <= SharedReg11_out;
SharedReg10_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_43_cast <= SharedReg10_out;
SharedReg9_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_44_cast <= SharedReg9_out;
SharedReg13_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_45_cast <= SharedReg13_out;
SharedReg809_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_46_cast <= SharedReg809_out;
SharedReg416_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_47_cast <= SharedReg416_out;
SharedReg146_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_48_cast <= SharedReg146_out;
SharedReg671_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_49_cast <= SharedReg671_out;
SharedReg4_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_50_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_51_cast <= SharedReg7_out;
SharedReg818_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_52_cast <= SharedReg818_out;
SharedReg410_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_53_cast <= SharedReg410_out;
SharedReg410_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_54_cast <= SharedReg410_out;
SharedReg431_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_55_cast <= SharedReg431_out;
SharedReg524_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_56_cast <= SharedReg524_out;
SharedReg874_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_57_cast <= SharedReg874_out;
SharedReg677_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_58_cast <= SharedReg677_out;
SharedReg549_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_59_cast <= SharedReg549_out;
Delay43No5_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_60_cast <= Delay43No5_out;
SharedReg313_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_61_cast <= SharedReg313_out;
SharedReg519_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_62_cast <= SharedReg519_out;
SharedReg801_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_63_cast <= SharedReg801_out;
SharedReg819_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_64_cast <= SharedReg819_out;
   MUX_Add2_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg410_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg521_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg416_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg685_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg830_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg174_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg410_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg140_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg410_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg302_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg417_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg519_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg663_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg859_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg519_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg425_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg807_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg142_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg808_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg312_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg872_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg937_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg292_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg312_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg146_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg865_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg806_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg424_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg412_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg412_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg803_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg2_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg17_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg425_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg695_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg11_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg10_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg9_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg13_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg809_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg416_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg146_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg671_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg4_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg672_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg7_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg818_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg410_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg410_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg431_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg524_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg874_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg677_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg549_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => Delay43No5_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg150_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg313_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg519_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg801_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg819_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg150_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg425_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg534_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add2_4_impl_0_out);

   Delay1No40_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_4_impl_0_out,
                 Y => Delay1No40_out);

SharedReg805_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg805_out;
SharedReg801_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg801_out;
SharedReg703_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg703_out;
SharedReg184_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg184_out;
SharedReg536_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg536_out;
SharedReg661_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg661_out;
SharedReg139_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg139_out;
SharedReg286_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg286_out;
SharedReg541_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg541_out;
SharedReg806_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg806_out;
SharedReg414_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg414_out;
SharedReg690_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg690_out;
SharedReg820_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg820_out;
SharedReg139_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg139_out;
SharedReg803_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg803_out;
SharedReg158_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg158_out;
SharedReg520_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg520_out;
SharedReg139_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg139_out;
SharedReg410_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg410_out;
SharedReg809_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg809_out;
SharedReg702_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg702_out;
SharedReg801_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg801_out;
SharedReg536_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg536_out;
SharedReg801_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg801_out;
SharedReg139_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg139_out;
SharedReg411_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg411_out;
SharedReg328_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg328_out;
SharedReg711_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg711_out;
SharedReg855_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_29_cast <= SharedReg855_out;
SharedReg140_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_30_cast <= SharedReg140_out;
SharedReg139_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_31_cast <= SharedReg139_out;
SharedReg856_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_32_cast <= SharedReg856_out;
SharedReg808_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_33_cast <= SharedReg808_out;
SharedReg523_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_34_cast <= SharedReg523_out;
SharedReg519_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_35_cast <= SharedReg519_out;
SharedReg519_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_36_cast <= SharedReg519_out;
SharedReg802_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_37_cast <= SharedReg802_out;
SharedReg18_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_38_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_39_cast <= SharedReg20_out;
SharedReg35_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_40_cast <= SharedReg35_out;
SharedReg686_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_41_cast <= SharedReg686_out;
SharedReg29_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_42_cast <= SharedReg29_out;
SharedReg28_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_43_cast <= SharedReg28_out;
SharedReg27_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_44_cast <= SharedReg27_out;
SharedReg31_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_45_cast <= SharedReg31_out;
SharedReg527_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_46_cast <= SharedReg527_out;
SharedReg523_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_47_cast <= SharedReg523_out;
SharedReg147_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_48_cast <= SharedReg147_out;
SharedReg672_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_49_cast <= SharedReg672_out;
SharedReg22_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_50_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_51_cast <= SharedReg25_out;
SharedReg419_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_52_cast <= SharedReg419_out;
SharedReg519_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_53_cast <= SharedReg519_out;
SharedReg417_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_54_cast <= SharedReg417_out;
SharedReg542_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_55_cast <= SharedReg542_out;
SharedReg801_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_56_cast <= SharedReg801_out;
SharedReg857_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_57_cast <= SharedReg857_out;
SharedReg720_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_58_cast <= SharedReg720_out;
SharedReg832_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_59_cast <= SharedReg832_out;
SharedReg546_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_60_cast <= SharedReg546_out;
SharedReg308_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_61_cast <= SharedReg308_out;
SharedReg801_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_62_cast <= SharedReg801_out;
SharedReg523_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_63_cast <= SharedReg523_out;
SharedReg542_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_64_cast <= SharedReg542_out;
   MUX_Add2_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg805_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg801_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg414_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg690_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg820_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg139_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg803_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg158_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg520_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg139_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg410_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg809_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg703_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg702_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg801_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg536_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg801_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg139_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg411_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg328_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg711_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg855_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg140_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg184_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg139_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg856_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg808_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg523_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg519_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg519_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg802_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg18_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg20_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg35_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg536_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg686_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg29_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg28_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg27_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg31_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg527_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg523_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg147_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg672_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg22_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg661_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg25_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg419_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg519_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg417_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg542_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg801_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg857_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg720_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg832_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg546_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg139_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg308_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg801_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg523_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg542_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg286_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg541_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg806_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add2_4_impl_1_out);

   Delay1No41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_4_impl_1_out,
                 Y => Delay1No41_out);

Delay1No42_out_to_Add2_5_impl_parent_implementedSystem_port_0_cast <= Delay1No42_out;
Delay1No43_out_to_Add2_5_impl_parent_implementedSystem_port_1_cast <= Delay1No43_out;
   Add2_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_5_impl_out,
                 X => Delay1No42_out_to_Add2_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No43_out_to_Add2_5_impl_parent_implementedSystem_port_1_cast);

SharedReg_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg_out;
SharedReg2_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg2_out;
SharedReg2_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg2_out;
SharedReg8_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg8_out;
SharedReg9_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg9_out;
SharedReg10_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg10_out;
SharedReg13_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg13_out;
SharedReg15_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg15_out;
SharedReg17_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg17_out;
SharedReg17_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg17_out;
SharedReg721_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg721_out;
SharedReg321_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg321_out;
SharedReg696_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg696_out;
SharedReg321_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_14_cast <= SharedReg321_out;
SharedReg332_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_15_cast <= SharedReg332_out;
SharedReg535_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_16_cast <= SharedReg535_out;
SharedReg540_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_17_cast <= SharedReg540_out;
SharedReg440_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_18_cast <= SharedReg440_out;
SharedReg195_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_19_cast <= SharedReg195_out;
SharedReg425_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_20_cast <= SharedReg425_out;
SharedReg695_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_21_cast <= SharedReg695_out;
SharedReg202_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_22_cast <= SharedReg202_out;
SharedReg340_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_23_cast <= SharedReg340_out;
SharedReg439_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_24_cast <= SharedReg439_out;
SharedReg993_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_25_cast <= SharedReg993_out;
SharedReg168_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_26_cast <= SharedReg168_out;
SharedReg425_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_27_cast <= SharedReg425_out;
SharedReg826_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_28_cast <= SharedReg826_out;
SharedReg535_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_29_cast <= SharedReg535_out;
SharedReg551_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_30_cast <= SharedReg551_out;
SharedReg700_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_31_cast <= SharedReg700_out;
SharedReg316_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_32_cast <= SharedReg316_out;
SharedReg861_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_33_cast <= SharedReg861_out;
SharedReg565_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_34_cast <= SharedReg565_out;
SharedReg166_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_35_cast <= SharedReg166_out;
SharedReg825_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_36_cast <= SharedReg825_out;
SharedReg425_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_37_cast <= SharedReg425_out;
SharedReg884_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_38_cast <= SharedReg884_out;
SharedReg535_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_39_cast <= SharedReg535_out;
SharedReg334_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_40_cast <= SharedReg334_out;
SharedReg433_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_41_cast <= SharedReg433_out;
SharedReg167_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_42_cast <= SharedReg167_out;
SharedReg828_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_43_cast <= SharedReg828_out;
SharedReg846_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_44_cast <= SharedReg846_out;
SharedReg825_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_45_cast <= SharedReg825_out;
SharedReg541_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_46_cast <= SharedReg541_out;
SharedReg164_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_47_cast <= SharedReg164_out;
SharedReg550_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_48_cast <= SharedReg550_out;
SharedReg427_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_49_cast <= SharedReg427_out;
SharedReg448_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_50_cast <= SharedReg448_out;
SharedReg188_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_51_cast <= SharedReg188_out;
SharedReg188_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_52_cast <= SharedReg188_out;
SharedReg883_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_53_cast <= SharedReg883_out;
SharedReg337_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_54_cast <= SharedReg337_out;
SharedReg431_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_55_cast <= SharedReg431_out;
SharedReg427_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_56_cast <= SharedReg427_out;
SharedReg442_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_57_cast <= SharedReg442_out;
SharedReg689_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_58_cast <= SharedReg689_out;
SharedReg821_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_59_cast <= SharedReg821_out;
SharedReg537_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_60_cast <= SharedReg537_out;
SharedReg848_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_61_cast <= SharedReg848_out;
SharedReg823_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_62_cast <= SharedReg823_out;
SharedReg819_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_63_cast <= SharedReg819_out;
   MUX_Add2_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_63_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg2_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg721_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg321_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg696_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg321_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg332_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg535_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg540_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg440_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg195_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg425_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg2_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg695_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg202_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg340_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg439_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg993_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg168_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg425_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg826_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg535_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg551_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg8_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg700_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg316_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg861_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg565_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg166_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg825_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg425_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg884_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg535_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg334_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg9_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg433_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg167_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg828_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg846_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg825_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg541_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg164_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg550_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg427_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg448_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg10_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg188_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg188_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg883_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg337_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg431_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg427_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg442_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg689_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg821_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg537_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg13_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg848_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg823_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg819_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_63_cast,
                 iS_7 => SharedReg15_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg17_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg17_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Add2_5_impl_0_LUT_out,
                 oMux => MUX_Add2_5_impl_0_out);

   Delay1No42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_5_impl_0_out,
                 Y => Delay1No42_out);

SharedReg18_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg20_out;
SharedReg20_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg20_out;
SharedReg26_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg26_out;
SharedReg27_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg27_out;
SharedReg28_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg28_out;
SharedReg31_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg31_out;
SharedReg33_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg33_out;
SharedReg35_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg35_out;
SharedReg35_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg35_out;
SharedReg819_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg819_out;
SharedReg338_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg338_out;
SharedReg819_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg819_out;
SharedReg553_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_14_cast <= SharedReg553_out;
SharedReg536_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_15_cast <= SharedReg536_out;
SharedReg539_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_16_cast <= SharedReg539_out;
SharedReg821_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_17_cast <= SharedReg821_out;
SharedReg687_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_18_cast <= SharedReg687_out;
SharedReg850_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_19_cast <= SharedReg850_out;
SharedReg663_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_20_cast <= SharedReg663_out;
SharedReg332_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_21_cast <= SharedReg332_out;
SharedReg426_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_22_cast <= SharedReg426_out;
SharedReg708_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_23_cast <= SharedReg708_out;
SharedReg819_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_24_cast <= SharedReg819_out;
SharedReg837_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_25_cast <= SharedReg837_out;
SharedReg164_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_26_cast <= SharedReg164_out;
SharedReg819_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_27_cast <= SharedReg819_out;
SharedReg685_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_28_cast <= SharedReg685_out;
SharedReg823_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_29_cast <= SharedReg823_out;
SharedReg341_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_30_cast <= SharedReg341_out;
SharedReg994_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_31_cast <= SharedReg994_out;
SharedReg163_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_32_cast <= SharedReg163_out;
SharedReg827_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_33_cast <= SharedReg827_out;
SharedReg206_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_34_cast <= SharedReg206_out;
SharedReg836_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_35_cast <= SharedReg836_out;
SharedReg162_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_36_cast <= SharedReg162_out;
SharedReg544_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_37_cast <= SharedReg544_out;
SharedReg560_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_38_cast <= SharedReg560_out;
SharedReg349_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_39_cast <= SharedReg349_out;
SharedReg827_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_40_cast <= SharedReg827_out;
SharedReg824_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_41_cast <= SharedReg824_out;
SharedReg181_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_42_cast <= SharedReg181_out;
SharedReg824_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_43_cast <= SharedReg824_out;
SharedReg535_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_44_cast <= SharedReg535_out;
SharedReg311_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_45_cast <= SharedReg311_out;
SharedReg440_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_46_cast <= SharedReg440_out;
SharedReg707_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_47_cast <= SharedReg707_out;
SharedReg206_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_48_cast <= SharedReg206_out;
SharedReg344_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_49_cast <= SharedReg344_out;
SharedReg899_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_50_cast <= SharedReg899_out;
SharedReg429_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_51_cast <= SharedReg429_out;
SharedReg183_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_52_cast <= SharedReg183_out;
SharedReg903_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_53_cast <= SharedReg903_out;
SharedReg535_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_54_cast <= SharedReg535_out;
SharedReg551_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_55_cast <= SharedReg551_out;
SharedReg820_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_56_cast <= SharedReg820_out;
SharedReg163_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_57_cast <= SharedReg163_out;
SharedReg819_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_58_cast <= SharedReg819_out;
SharedReg163_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_59_cast <= SharedReg163_out;
SharedReg838_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_60_cast <= SharedReg838_out;
SharedReg539_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_61_cast <= SharedReg539_out;
SharedReg711_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_62_cast <= SharedReg711_out;
SharedReg535_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_63_cast <= SharedReg535_out;
   MUX_Add2_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_63_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg18_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg20_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg819_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg338_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg819_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg553_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg536_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg539_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg821_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg687_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg850_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg663_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg20_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg332_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg426_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg708_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg819_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg837_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg164_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg819_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg685_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg823_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg341_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg26_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg994_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg163_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg827_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg206_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg836_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg162_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg544_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg560_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg349_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg827_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg27_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg824_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg181_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg824_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg535_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg311_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg440_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg707_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg206_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg344_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg899_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg28_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg429_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg183_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg903_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg535_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg551_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg820_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg163_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg819_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg163_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg838_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg31_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg539_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg711_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg535_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_63_cast,
                 iS_7 => SharedReg33_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg35_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg35_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Add2_5_impl_1_LUT_out,
                 oMux => MUX_Add2_5_impl_1_out);

   Delay1No43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_5_impl_1_out,
                 Y => Delay1No43_out);

Delay1No44_out_to_Add2_6_impl_parent_implementedSystem_port_0_cast <= Delay1No44_out;
Delay1No45_out_to_Add2_6_impl_parent_implementedSystem_port_1_cast <= Delay1No45_out;
   Add2_6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_6_impl_out,
                 X => Delay1No44_out_to_Add2_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No45_out_to_Add2_6_impl_parent_implementedSystem_port_1_cast);

SharedReg_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg_out;
SharedReg1_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1_out;
SharedReg3_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg3_out;
SharedReg3_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg3_out;
SharedReg7_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg7_out;
SharedReg8_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg8_out;
SharedReg9_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg9_out;
SharedReg10_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg10_out;
SharedReg12_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg12_out;
SharedReg16_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg16_out;
SharedReg321_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg321_out;
SharedReg440_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg440_out;
SharedReg891_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_13_cast <= SharedReg891_out;
SharedReg203_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_14_cast <= SharedReg203_out;
SharedReg446_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_15_cast <= SharedReg446_out;
SharedReg894_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_16_cast <= SharedReg894_out;
SharedReg440_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_17_cast <= SharedReg440_out;
SharedReg454_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_18_cast <= SharedReg454_out;
SharedReg177_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_19_cast <= SharedReg177_out;
SharedReg191_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_20_cast <= SharedReg191_out;
SharedReg440_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_21_cast <= SharedReg440_out;
SharedReg191_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_22_cast <= SharedReg191_out;
SharedReg451_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_23_cast <= SharedReg451_out;
SharedReg440_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_24_cast <= SharedReg440_out;
SharedReg888_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_25_cast <= SharedReg888_out;
SharedReg553_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_26_cast <= SharedReg553_out;
SharedReg898_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_27_cast <= SharedReg898_out;
SharedReg888_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_28_cast <= SharedReg888_out;
SharedReg179_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_29_cast <= SharedReg179_out;
SharedReg700_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_30_cast <= SharedReg700_out;
SharedReg193_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_31_cast <= SharedReg193_out;
SharedReg440_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_32_cast <= SharedReg440_out;
SharedReg332_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_33_cast <= SharedReg332_out;
SharedReg446_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_34_cast <= SharedReg446_out;
SharedReg885_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_35_cast <= SharedReg885_out;
SharedReg446_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_36_cast <= SharedReg446_out;
SharedReg987_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_37_cast <= SharedReg987_out;
SharedReg883_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_38_cast <= SharedReg883_out;
SharedReg843_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_39_cast <= SharedReg843_out;
SharedReg854_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_40_cast <= SharedReg854_out;
SharedReg557_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_41_cast <= SharedReg557_out;
SharedReg987_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_42_cast <= SharedReg987_out;
SharedReg987_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_43_cast <= SharedReg987_out;
SharedReg555_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_44_cast <= SharedReg555_out;
SharedReg886_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_45_cast <= SharedReg886_out;
SharedReg553_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_46_cast <= SharedReg553_out;
SharedReg837_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_47_cast <= SharedReg837_out;
SharedReg337_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_48_cast <= SharedReg337_out;
   MUX_Add2_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_48_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg321_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg440_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg891_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg203_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg446_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg894_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg440_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg454_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg177_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg191_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg3_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg440_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg191_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg451_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg440_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg888_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg553_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg898_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg888_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg179_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg700_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg3_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg193_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg440_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg332_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg446_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg885_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg446_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg987_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg883_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg843_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg854_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg7_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg557_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg987_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg987_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg555_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg886_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg553_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg837_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg337_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_48_cast,
                 iS_5 => SharedReg8_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg9_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg10_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg12_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg16_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Add2_6_impl_0_LUT_out,
                 oMux => MUX_Add2_6_impl_0_out);

   Delay1No44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_6_impl_0_out,
                 Y => Delay1No44_out);

SharedReg25_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg25_out;
SharedReg18_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg18_out;
SharedReg19_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg19_out;
SharedReg21_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg21_out;
SharedReg21_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg21_out;
SharedReg26_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg26_out;
SharedReg27_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg27_out;
SharedReg28_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg28_out;
SharedReg30_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg30_out;
SharedReg34_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg34_out;
SharedReg551_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg551_out;
SharedReg551_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg551_out;
SharedReg332_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_13_cast <= SharedReg332_out;
SharedReg886_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_14_cast <= SharedReg886_out;
SharedReg557_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_15_cast <= SharedReg557_out;
SharedReg186_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_16_cast <= SharedReg186_out;
SharedReg447_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_17_cast <= SharedReg447_out;
SharedReg685_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_18_cast <= SharedReg685_out;
SharedReg552_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_19_cast <= SharedReg552_out;
SharedReg551_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_20_cast <= SharedReg551_out;
SharedReg336_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_21_cast <= SharedReg336_out;
SharedReg552_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_22_cast <= SharedReg552_out;
SharedReg837_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_23_cast <= SharedReg837_out;
SharedReg332_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_24_cast <= SharedReg332_out;
SharedReg882_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_25_cast <= SharedReg882_out;
SharedReg310_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_26_cast <= SharedReg310_out;
SharedReg709_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_27_cast <= SharedReg709_out;
SharedReg839_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_28_cast <= SharedReg839_out;
SharedReg168_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_29_cast <= SharedReg168_out;
SharedReg333_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_30_cast <= SharedReg333_out;
SharedReg984_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_31_cast <= SharedReg984_out;
SharedReg555_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_32_cast <= SharedReg555_out;
SharedReg558_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_33_cast <= SharedReg558_out;
SharedReg905_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_34_cast <= SharedReg905_out;
SharedReg1002_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_35_cast <= SharedReg1002_out;
SharedReg842_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_36_cast <= SharedReg842_out;
SharedReg900_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_37_cast <= SharedReg900_out;
SharedReg164_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_38_cast <= SharedReg164_out;
SharedReg449_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_39_cast <= SharedReg449_out;
SharedReg842_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_40_cast <= SharedReg842_out;
SharedReg1000_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_41_cast <= SharedReg1000_out;
SharedReg188_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_42_cast <= SharedReg188_out;
SharedReg903_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_43_cast <= SharedReg903_out;
SharedReg841_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_44_cast <= SharedReg841_out;
SharedReg987_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_45_cast <= SharedReg987_out;
SharedReg837_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_46_cast <= SharedReg837_out;
SharedReg707_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_47_cast <= SharedReg707_out;
SharedReg555_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_48_cast <= SharedReg555_out;
   MUX_Add2_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_48_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg25_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg18_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg551_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg551_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg332_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg886_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg557_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg186_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg447_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg685_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg552_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg551_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg19_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg336_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg552_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg837_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg332_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg882_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg310_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg709_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg839_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg168_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg333_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg21_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg984_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg555_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg558_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg905_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1002_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg842_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg900_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg164_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg449_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg842_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg21_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1000_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg188_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg903_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg841_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg987_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg837_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg707_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg555_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_48_cast,
                 iS_5 => SharedReg26_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg27_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg28_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg30_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg34_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Add2_6_impl_1_LUT_out,
                 oMux => MUX_Add2_6_impl_1_out);

   Delay1No45_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_6_impl_1_out,
                 Y => Delay1No45_out);

Delay1No46_out_to_Add11_0_impl_parent_implementedSystem_port_0_cast <= Delay1No46_out;
Delay1No47_out_to_Add11_0_impl_parent_implementedSystem_port_1_cast <= Delay1No47_out;
   Add11_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_0_impl_out,
                 X => Delay1No46_out_to_Add11_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No47_out_to_Add11_0_impl_parent_implementedSystem_port_1_cast);

SharedReg731_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg731_out;
SharedReg1_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1_out;
SharedReg3_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg3_out;
SharedReg17_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg17_out;
SharedReg15_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg15_out;
SharedReg11_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg11_out;
SharedReg12_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg12_out;
SharedReg16_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg16_out;
SharedReg8_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg8_out;
SharedReg737_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg737_out;
SharedReg461_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg461_out;
SharedReg735_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg735_out;
SharedReg576_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg576_out;
SharedReg469_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg469_out;
Delay43No_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_15_cast <= Delay43No_out;
SharedReg733_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg733_out;
SharedReg358_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg358_out;
SharedReg738_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg738_out;
SharedReg729_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg729_out;
SharedReg460_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg460_out;
SharedReg586_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg586_out;
SharedReg210_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg210_out;
SharedReg38_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg38_out;
SharedReg350_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg350_out;
SharedReg211_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg211_out;
SharedReg455_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg455_out;
SharedReg729_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg729_out;
SharedReg225_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg225_out;
SharedReg350_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_29_cast <= SharedReg350_out;
SharedReg457_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_30_cast <= SharedReg457_out;
SharedReg208_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_31_cast <= SharedReg208_out;
SharedReg740_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_32_cast <= SharedReg740_out;
SharedReg220_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_33_cast <= SharedReg220_out;
SharedReg577_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_34_cast <= SharedReg577_out;
SharedReg49_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_35_cast <= SharedReg49_out;
SharedReg49_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_36_cast <= SharedReg49_out;
SharedReg579_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_37_cast <= SharedReg579_out;
SharedReg470_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_38_cast <= SharedReg470_out;
SharedReg356_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_39_cast <= SharedReg356_out;
SharedReg593_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_40_cast <= SharedReg593_out;
SharedReg758_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_41_cast <= SharedReg758_out;
SharedReg910_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_42_cast <= SharedReg910_out;
SharedReg350_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_43_cast <= SharedReg350_out;
SharedReg209_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_44_cast <= SharedReg209_out;
SharedReg350_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_45_cast <= SharedReg350_out;
SharedReg350_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_46_cast <= SharedReg350_out;
SharedReg357_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_47_cast <= SharedReg357_out;
SharedReg455_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_48_cast <= SharedReg455_out;
SharedReg571_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_49_cast <= SharedReg571_out;
SharedReg455_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_50_cast <= SharedReg455_out;
SharedReg365_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_51_cast <= SharedReg365_out;
SharedReg735_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_52_cast <= SharedReg735_out;
SharedReg213_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_53_cast <= SharedReg213_out;
SharedReg736_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_54_cast <= SharedReg736_out;
SharedReg64_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_55_cast <= SharedReg64_out;
SharedReg610_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_56_cast <= SharedReg610_out;
SharedReg910_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_57_cast <= SharedReg910_out;
SharedReg239_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_58_cast <= SharedReg239_out;
SharedReg67_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_59_cast <= SharedReg67_out;
SharedReg365_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_60_cast <= SharedReg365_out;
SharedReg213_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_61_cast <= SharedReg213_out;
SharedReg963_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_62_cast <= SharedReg963_out;
SharedReg599_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_63_cast <= SharedReg599_out;
SharedReg376_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_64_cast <= SharedReg376_out;
   MUX_Add11_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg731_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg461_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg735_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg576_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg469_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => Delay43No_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg733_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg358_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg738_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg729_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg460_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg3_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg586_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg210_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg38_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg350_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg211_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg455_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg729_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg225_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg350_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg457_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg17_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg208_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg740_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg220_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg577_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg49_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg49_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg579_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg470_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg356_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg593_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg15_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg758_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg910_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg350_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg209_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg350_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg350_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg357_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg455_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg571_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg455_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg11_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg365_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg735_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg213_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg736_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg64_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg610_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg910_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg239_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg67_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg365_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg12_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg213_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg963_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg599_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg376_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg16_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg8_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg737_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add11_0_impl_0_out);

   Delay1No46_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_0_impl_0_out,
                 Y => Delay1No46_out);

SharedReg730_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg730_out;
SharedReg19_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg19_out;
SharedReg21_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg21_out;
SharedReg35_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg35_out;
SharedReg33_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg33_out;
SharedReg29_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg30_out;
SharedReg34_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg34_out;
SharedReg26_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg26_out;
SharedReg463_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg463_out;
SharedReg737_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg737_out;
SharedReg734_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg734_out;
SharedReg577_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg577_out;
SharedReg742_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg742_out;
SharedReg466_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg466_out;
SharedReg455_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg455_out;
SharedReg746_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg746_out;
SharedReg464_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg464_out;
SharedReg462_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg462_out;
SharedReg729_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg729_out;
SharedReg959_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg959_out;
SharedReg60_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg60_out;
SharedReg232_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg232_out;
SharedReg456_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg456_out;
SharedReg61_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg61_out;
SharedReg729_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg729_out;
SharedReg459_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg459_out;
SharedReg62_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg62_out;
SharedReg733_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_29_cast <= SharedReg733_out;
SharedReg729_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_30_cast <= SharedReg729_out;
SharedReg214_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_31_cast <= SharedReg214_out;
SharedReg730_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_32_cast <= SharedReg730_out;
SharedReg36_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_33_cast <= SharedReg36_out;
SharedReg957_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_34_cast <= SharedReg957_out;
SharedReg208_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_35_cast <= SharedReg208_out;
SharedReg37_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_36_cast <= SharedReg37_out;
SharedReg567_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_37_cast <= SharedReg567_out;
SharedReg734_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_38_cast <= SharedReg734_out;
SharedReg354_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_39_cast <= SharedReg354_out;
SharedReg598_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_40_cast <= SharedReg598_out;
SharedReg748_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_41_cast <= SharedReg748_out;
SharedReg597_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_42_cast <= SharedReg597_out;
SharedReg731_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_43_cast <= SharedReg731_out;
SharedReg57_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_44_cast <= SharedReg57_out;
SharedReg456_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_45_cast <= SharedReg456_out;
SharedReg731_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_46_cast <= SharedReg731_out;
SharedReg350_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_47_cast <= SharedReg350_out;
SharedReg737_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_48_cast <= SharedReg737_out;
SharedReg980_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_49_cast <= SharedReg980_out;
SharedReg729_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_50_cast <= SharedReg729_out;
SharedReg472_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_51_cast <= SharedReg472_out;
SharedReg729_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_52_cast <= SharedReg729_out;
SharedReg208_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_53_cast <= SharedReg208_out;
SharedReg351_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_54_cast <= SharedReg351_out;
SharedReg253_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_55_cast <= SharedReg253_out;
SharedReg910_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_56_cast <= SharedReg910_out;
SharedReg614_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_57_cast <= SharedReg614_out;
SharedReg85_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_58_cast <= SharedReg85_out;
SharedReg256_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_59_cast <= SharedReg256_out;
SharedReg473_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_60_cast <= SharedReg473_out;
SharedReg62_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_61_cast <= SharedReg62_out;
SharedReg957_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_62_cast <= SharedReg957_out;
SharedReg594_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_63_cast <= SharedReg594_out;
SharedReg471_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_64_cast <= SharedReg471_out;
   MUX_Add11_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg730_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg19_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg737_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg734_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg577_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg742_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg466_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg455_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg746_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg464_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg462_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg729_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg21_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg959_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg60_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg232_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg456_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg61_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg729_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg459_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg62_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg733_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg729_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg35_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg214_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg730_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg36_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg957_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg208_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg37_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg567_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg734_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg354_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg598_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg33_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg748_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg597_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg731_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg57_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg456_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg731_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg350_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg737_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg980_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg729_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg29_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg472_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg729_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg208_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg351_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg253_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg910_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg614_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg85_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg256_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg473_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg30_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg62_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg957_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg594_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg471_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg34_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg26_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg463_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add11_0_impl_1_out);

   Delay1No47_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_0_impl_1_out,
                 Y => Delay1No47_out);

Delay1No48_out_to_Add11_1_impl_parent_implementedSystem_port_0_cast <= Delay1No48_out;
Delay1No49_out_to_Add11_1_impl_parent_implementedSystem_port_1_cast <= Delay1No49_out;
   Add11_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_1_impl_out,
                 X => Delay1No48_out_to_Add11_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No49_out_to_Add11_1_impl_parent_implementedSystem_port_1_cast);

SharedReg635_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg635_out;
SharedReg621_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg621_out;
SharedReg92_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg92_out;
SharedReg239_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg239_out;
SharedReg380_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg380_out;
SharedReg67_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg67_out;
SharedReg599_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg599_out;
SharedReg912_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg912_out;
SharedReg391_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg391_out;
SharedReg749_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg749_out;
SharedReg1_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1_out;
SharedReg3_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg3_out;
SharedReg17_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg17_out;
SharedReg15_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg15_out;
SharedReg11_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg11_out;
SharedReg12_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg12_out;
SharedReg16_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg16_out;
SharedReg8_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg8_out;
SharedReg755_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg755_out;
SharedReg477_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg477_out;
SharedReg753_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg753_out;
SharedReg602_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg602_out;
SharedReg485_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg485_out;
Delay43No1_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_24_cast <= Delay43No1_out;
SharedReg751_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg751_out;
SharedReg373_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg373_out;
SharedReg756_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg756_out;
SharedReg386_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg386_out;
SharedReg476_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_29_cast <= SharedReg476_out;
SharedReg975_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_30_cast <= SharedReg975_out;
SharedReg236_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_31_cast <= SharedReg236_out;
SharedReg64_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_32_cast <= SharedReg64_out;
SharedReg365_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_33_cast <= SharedReg365_out;
SharedReg237_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_34_cast <= SharedReg237_out;
SharedReg471_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_35_cast <= SharedReg471_out;
SharedReg747_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_36_cast <= SharedReg747_out;
SharedReg251_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_37_cast <= SharedReg251_out;
SharedReg365_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_38_cast <= SharedReg365_out;
SharedReg473_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_39_cast <= SharedReg473_out;
SharedReg933_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_40_cast <= SharedReg933_out;
SharedReg90_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_41_cast <= SharedReg90_out;
SharedReg108_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_42_cast <= SharedReg108_out;
SharedReg603_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_43_cast <= SharedReg603_out;
SharedReg75_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_44_cast <= SharedReg75_out;
SharedReg75_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_45_cast <= SharedReg75_out;
SharedReg605_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_46_cast <= SharedReg605_out;
SharedReg486_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_47_cast <= SharedReg486_out;
SharedReg371_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_48_cast <= SharedReg371_out;
SharedReg617_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_49_cast <= SharedReg617_out;
SharedReg776_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_50_cast <= SharedReg776_out;
SharedReg272_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_51_cast <= SharedReg272_out;
SharedReg365_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_52_cast <= SharedReg365_out;
SharedReg235_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_53_cast <= SharedReg235_out;
SharedReg365_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_54_cast <= SharedReg365_out;
SharedReg103_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_55_cast <= SharedReg103_out;
SharedReg394_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_56_cast <= SharedReg394_out;
SharedReg493_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_57_cast <= SharedReg493_out;
SharedReg491_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_58_cast <= SharedReg491_out;
SharedReg866_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_59_cast <= SharedReg866_out;
SharedReg935_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_60_cast <= SharedReg935_out;
SharedReg104_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_61_cast <= SharedReg104_out;
SharedReg907_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_62_cast <= SharedReg907_out;
SharedReg907_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_63_cast <= SharedReg907_out;
SharedReg380_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_64_cast <= SharedReg380_out;
   MUX_Add11_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg635_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg621_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg3_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg17_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg15_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg11_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg12_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg16_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg8_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg755_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg477_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg92_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg753_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg602_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg485_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => Delay43No1_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg751_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg373_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg756_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg386_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg476_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg975_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg239_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg236_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg64_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg365_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg237_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg471_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg747_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg251_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg365_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg473_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg933_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg380_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg90_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg108_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg603_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg75_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg75_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg605_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg486_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg371_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg617_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg776_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg67_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg272_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg365_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg235_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg365_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg103_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg394_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg493_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg491_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg866_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg935_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg599_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg104_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg907_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg907_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg380_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg912_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg391_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg749_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add11_1_impl_0_out);

   Delay1No48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_1_impl_0_out,
                 Y => Delay1No48_out);

SharedReg621_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg621_out;
SharedReg928_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg928_out;
SharedReg112_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg112_out;
SharedReg281_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg281_out;
SharedReg489_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg489_out;
SharedReg88_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg88_out;
SharedReg906_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg906_out;
SharedReg618_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg618_out;
SharedReg487_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg487_out;
SharedReg748_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg748_out;
SharedReg19_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg19_out;
SharedReg21_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg21_out;
SharedReg35_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg35_out;
SharedReg33_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg33_out;
SharedReg29_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg30_out;
SharedReg34_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg34_out;
SharedReg26_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg26_out;
SharedReg479_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg479_out;
SharedReg755_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg755_out;
SharedReg752_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg752_out;
SharedReg603_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg603_out;
SharedReg760_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg760_out;
SharedReg482_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg482_out;
SharedReg471_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg471_out;
SharedReg764_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg764_out;
SharedReg480_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg480_out;
SharedReg494_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg494_out;
SharedReg747_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_29_cast <= SharedReg747_out;
SharedReg908_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_30_cast <= SharedReg908_out;
SharedReg86_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_31_cast <= SharedReg86_out;
SharedReg257_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_32_cast <= SharedReg257_out;
SharedReg472_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_33_cast <= SharedReg472_out;
SharedReg87_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_34_cast <= SharedReg87_out;
SharedReg747_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_35_cast <= SharedReg747_out;
SharedReg475_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_36_cast <= SharedReg475_out;
SharedReg88_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_37_cast <= SharedReg88_out;
SharedReg751_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_38_cast <= SharedReg751_out;
SharedReg747_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_39_cast <= SharedReg747_out;
SharedReg638_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_40_cast <= SharedReg638_out;
SharedReg282_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_41_cast <= SharedReg282_out;
SharedReg265_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_42_cast <= SharedReg265_out;
SharedReg906_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_43_cast <= SharedReg906_out;
SharedReg234_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_44_cast <= SharedReg234_out;
SharedReg63_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_45_cast <= SharedReg63_out;
SharedReg567_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_46_cast <= SharedReg567_out;
SharedReg752_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_47_cast <= SharedReg752_out;
SharedReg369_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_48_cast <= SharedReg369_out;
SharedReg622_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_49_cast <= SharedReg622_out;
SharedReg766_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_50_cast <= SharedReg766_out;
SharedReg88_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_51_cast <= SharedReg88_out;
SharedReg749_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_52_cast <= SharedReg749_out;
SharedReg83_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_53_cast <= SharedReg83_out;
SharedReg472_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_54_cast <= SharedReg472_out;
SharedReg234_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_55_cast <= SharedReg234_out;
SharedReg387_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_56_cast <= SharedReg387_out;
SharedReg770_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_57_cast <= SharedReg770_out;
SharedReg769_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_58_cast <= SharedReg769_out;
SharedReg640_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_59_cast <= SharedReg640_out;
SharedReg621_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_60_cast <= SharedReg621_out;
SharedReg234_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_61_cast <= SharedReg234_out;
SharedReg637_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_62_cast <= SharedReg637_out;
SharedReg636_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_63_cast <= SharedReg636_out;
SharedReg767_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_64_cast <= SharedReg767_out;
   MUX_Add11_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg621_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg928_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg19_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg21_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg35_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg33_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg29_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg30_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg34_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg26_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg479_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg755_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg112_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg752_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg603_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg760_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg482_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg471_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg764_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg480_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg494_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg747_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg908_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg281_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg86_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg257_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg472_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg87_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg747_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg475_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg88_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg751_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg747_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg638_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg489_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg282_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg265_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg906_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg234_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg63_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg567_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg752_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg369_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg622_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg766_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg88_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg88_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg749_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg83_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg472_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg234_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg387_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg770_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg769_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg640_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg621_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg906_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg234_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg637_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg636_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg767_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg618_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg487_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg748_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add11_1_impl_1_out);

   Delay1No49_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_1_impl_1_out,
                 Y => Delay1No49_out);

Delay1No50_out_to_Add11_2_impl_parent_implementedSystem_port_0_cast <= Delay1No50_out;
Delay1No51_out_to_Add11_2_impl_parent_implementedSystem_port_1_cast <= Delay1No51_out;
   Add11_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_2_impl_out,
                 X => Delay1No50_out_to_Add11_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No51_out_to_Add11_2_impl_parent_implementedSystem_port_1_cast);

SharedReg409_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg409_out;
SharedReg509_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg509_out;
SharedReg507_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg507_out;
SharedReg696_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg696_out;
SharedReg644_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg644_out;
SharedReg129_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg129_out;
SharedReg932_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg932_out;
SharedReg932_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg932_out;
SharedReg395_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg395_out;
SharedReg947_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg947_out;
SharedReg644_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg644_out;
SharedReg118_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg118_out;
SharedReg265_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg265_out;
SharedReg395_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg395_out;
SharedReg92_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg92_out;
SharedReg623_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg623_out;
SharedReg937_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg937_out;
SharedReg406_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg406_out;
SharedReg767_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg767_out;
SharedReg1_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1_out;
SharedReg3_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg3_out;
SharedReg17_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg17_out;
SharedReg15_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg15_out;
SharedReg11_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg11_out;
SharedReg12_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg12_out;
SharedReg16_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg16_out;
SharedReg8_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg8_out;
SharedReg265_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg265_out;
SharedReg493_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_29_cast <= SharedReg493_out;
SharedReg771_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_30_cast <= SharedReg771_out;
SharedReg627_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_31_cast <= SharedReg627_out;
SharedReg501_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_32_cast <= SharedReg501_out;
Delay43No2_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_33_cast <= Delay43No2_out;
SharedReg769_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_34_cast <= SharedReg769_out;
SharedReg388_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_35_cast <= SharedReg388_out;
SharedReg774_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_36_cast <= SharedReg774_out;
SharedReg401_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_37_cast <= SharedReg401_out;
SharedReg492_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_38_cast <= SharedReg492_out;
SharedReg923_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_39_cast <= SharedReg923_out;
SharedReg633_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_40_cast <= SharedReg633_out;
SharedReg517_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_41_cast <= SharedReg517_out;
SharedReg505_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_42_cast <= SharedReg505_out;
SharedReg263_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_43_cast <= SharedReg263_out;
SharedReg487_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_44_cast <= SharedReg487_out;
SharedReg765_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_45_cast <= SharedReg765_out;
SharedReg278_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_46_cast <= SharedReg278_out;
SharedReg380_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_47_cast <= SharedReg380_out;
SharedReg489_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_48_cast <= SharedReg489_out;
SharedReg642_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_49_cast <= SharedReg642_out;
SharedReg116_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_50_cast <= SharedReg116_out;
SharedReg395_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_51_cast <= SharedReg395_out;
SharedReg628_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_52_cast <= SharedReg628_out;
SharedReg100_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_53_cast <= SharedReg100_out;
SharedReg100_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_54_cast <= SharedReg100_out;
SharedReg395_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_55_cast <= SharedReg395_out;
SharedReg118_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_56_cast <= SharedReg118_out;
SharedReg403_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_57_cast <= SharedReg403_out;
SharedReg285_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_58_cast <= SharedReg285_out;
SharedReg663_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_59_cast <= SharedReg663_out;
SharedReg156_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_60_cast <= SharedReg156_out;
SharedReg114_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_61_cast <= SharedReg114_out;
SharedReg649_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_62_cast <= SharedReg649_out;
SharedReg933_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_63_cast <= SharedReg933_out;
SharedReg651_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_64_cast <= SharedReg651_out;
   MUX_Add11_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg409_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg509_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg644_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg118_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg265_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg395_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg92_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg623_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg937_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg406_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg767_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg507_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg3_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg17_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg15_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg11_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg12_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg16_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg8_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg265_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg493_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg771_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg696_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg627_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg501_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => Delay43No2_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg769_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg388_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg774_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg401_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg492_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg923_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg633_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg644_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg517_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg505_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg263_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg487_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg765_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg278_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg380_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg489_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg642_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg116_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg129_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg395_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg628_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg100_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg100_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg395_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg118_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg403_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg285_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg663_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg156_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg932_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg114_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg649_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg933_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg651_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg932_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg395_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg947_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add11_2_impl_0_out);

   Delay1No50_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_2_impl_0_out,
                 Y => Delay1No50_out);

SharedReg402_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg402_out;
SharedReg788_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg788_out;
SharedReg787_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg787_out;
SharedReg855_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg855_out;
SharedReg935_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg935_out;
SharedReg260_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg260_out;
SharedReg658_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg658_out;
SharedReg657_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg657_out;
SharedReg785_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg785_out;
SharedReg644_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg644_out;
SharedReg954_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg954_out;
SharedReg137_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg137_out;
SharedReg137_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg137_out;
SharedReg505_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg505_out;
SharedReg114_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg114_out;
SharedReg931_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg931_out;
SharedReg641_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg641_out;
SharedReg503_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg503_out;
SharedReg766_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg766_out;
SharedReg19_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg19_out;
SharedReg21_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg21_out;
SharedReg35_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg35_out;
SharedReg33_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg33_out;
SharedReg29_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg30_out;
SharedReg34_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg34_out;
SharedReg26_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg26_out;
SharedReg117_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg117_out;
SharedReg773_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_29_cast <= SharedReg773_out;
SharedReg770_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_30_cast <= SharedReg770_out;
SharedReg628_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_31_cast <= SharedReg628_out;
SharedReg778_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_32_cast <= SharedReg778_out;
SharedReg498_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_33_cast <= SharedReg498_out;
SharedReg487_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_34_cast <= SharedReg487_out;
SharedReg782_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_35_cast <= SharedReg782_out;
SharedReg496_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_36_cast <= SharedReg496_out;
SharedReg510_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_37_cast <= SharedReg510_out;
SharedReg765_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_38_cast <= SharedReg765_out;
SharedReg933_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_39_cast <= SharedReg933_out;
SharedReg653_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_40_cast <= SharedReg653_out;
SharedReg796_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_41_cast <= SharedReg796_out;
SharedReg783_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_42_cast <= SharedReg783_out;
SharedReg258_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_43_cast <= SharedReg258_out;
SharedReg765_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_44_cast <= SharedReg765_out;
SharedReg491_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_45_cast <= SharedReg491_out;
SharedReg88_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_46_cast <= SharedReg88_out;
SharedReg769_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_47_cast <= SharedReg769_out;
SharedReg765_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_48_cast <= SharedReg765_out;
SharedReg659_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_49_cast <= SharedReg659_out;
SharedReg307_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_50_cast <= SharedReg307_out;
SharedReg504_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_51_cast <= SharedReg504_out;
SharedReg931_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_52_cast <= SharedReg931_out;
SharedReg260_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_53_cast <= SharedReg260_out;
SharedReg89_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_54_cast <= SharedReg89_out;
SharedReg509_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_55_cast <= SharedReg509_out;
SharedReg260_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_56_cast <= SharedReg260_out;
SharedReg395_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_57_cast <= SharedReg395_out;
SharedReg291_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_58_cast <= SharedReg291_out;
SharedReg704_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_59_cast <= SharedReg704_out;
SharedReg290_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_60_cast <= SharedReg290_out;
SharedReg287_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_61_cast <= SharedReg287_out;
SharedReg931_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_62_cast <= SharedReg931_out;
SharedReg859_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_63_cast <= SharedReg859_out;
SharedReg906_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_64_cast <= SharedReg906_out;
   MUX_Add11_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg402_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg788_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg954_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg137_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg137_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg505_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg114_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg931_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg641_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg503_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg766_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg19_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg787_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg21_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg35_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg33_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg29_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg30_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg34_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg26_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg117_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg773_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg770_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg855_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg628_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg778_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg498_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg487_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg782_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg496_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg510_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg765_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg933_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg653_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg935_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg796_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg783_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg258_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg765_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg491_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg88_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg769_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg765_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg659_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg307_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg260_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg504_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg931_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg260_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg89_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg509_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg260_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg395_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg291_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg704_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg290_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg658_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg287_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg931_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg859_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg906_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg657_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg785_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg644_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add11_2_impl_1_out);

   Delay1No51_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_2_impl_1_out,
                 Y => Delay1No51_out);

Delay1No52_out_to_Add11_3_impl_parent_implementedSystem_port_0_cast <= Delay1No52_out;
Delay1No53_out_to_Add11_3_impl_parent_implementedSystem_port_1_cast <= Delay1No53_out;
   Add11_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_3_impl_out,
                 X => Delay1No52_out_to_Add11_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No53_out_to_Add11_3_impl_parent_implementedSystem_port_1_cast);

SharedReg290_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg290_out;
SharedReg418_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg418_out;
SharedReg139_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg139_out;
SharedReg687_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg687_out;
SharedReg179_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg179_out;
SharedReg139_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg139_out;
SharedReg865_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg865_out;
SharedReg857_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg857_out;
SharedReg868_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg868_out;
SharedReg424_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg424_out;
SharedReg525_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg525_out;
SharedReg523_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg523_out;
SharedReg717_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg717_out;
SharedReg665_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg665_out;
SharedReg303_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg303_out;
SharedReg856_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg856_out;
SharedReg856_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg856_out;
SharedReg410_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg410_out;
SharedReg656_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg656_out;
SharedReg665_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg665_out;
SharedReg142_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg142_out;
SharedReg290_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg290_out;
SharedReg410_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg410_out;
SharedReg118_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg118_out;
SharedReg646_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg646_out;
SharedReg861_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg861_out;
SharedReg421_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg421_out;
SharedReg410_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg410_out;
SharedReg1_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1_out;
SharedReg3_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_30_cast <= SharedReg3_out;
SharedReg17_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_31_cast <= SharedReg17_out;
SharedReg15_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_32_cast <= SharedReg15_out;
SharedReg11_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_33_cast <= SharedReg11_out;
SharedReg12_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_34_cast <= SharedReg12_out;
SharedReg16_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_35_cast <= SharedReg16_out;
SharedReg8_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_36_cast <= SharedReg8_out;
SharedReg290_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_37_cast <= SharedReg290_out;
SharedReg509_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_38_cast <= SharedReg509_out;
SharedReg789_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_39_cast <= SharedReg789_out;
SharedReg5_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_40_cast <= SharedReg5_out;
SharedReg15_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_41_cast <= SharedReg15_out;
SharedReg7_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_42_cast <= SharedReg7_out;
SharedReg787_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_43_cast <= SharedReg787_out;
SharedReg403_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_44_cast <= SharedReg403_out;
SharedReg792_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_45_cast <= SharedReg792_out;
SharedReg416_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_46_cast <= SharedReg416_out;
SharedReg508_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_47_cast <= SharedReg508_out;
SharedReg949_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_48_cast <= SharedReg949_out;
SharedReg654_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_49_cast <= SharedReg654_out;
SharedReg533_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_50_cast <= SharedReg533_out;
Delay43No4_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_51_cast <= Delay43No4_out;
SharedReg288_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_52_cast <= SharedReg288_out;
SharedReg503_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_53_cast <= SharedReg503_out;
SharedReg783_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_54_cast <= SharedReg783_out;
SharedReg801_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_55_cast <= SharedReg801_out;
SharedReg416_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_56_cast <= SharedReg416_out;
SharedReg873_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_57_cast <= SharedReg873_out;
SharedReg287_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_58_cast <= SharedReg287_out;
SharedReg546_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_59_cast <= SharedReg546_out;
SharedReg537_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_60_cast <= SharedReg537_out;
SharedReg664_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_61_cast <= SharedReg664_out;
SharedReg689_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_62_cast <= SharedReg689_out;
SharedReg314_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_63_cast <= SharedReg314_out;
SharedReg326_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_64_cast <= SharedReg326_out;
   MUX_Add11_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg290_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg418_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg525_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg523_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg717_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg665_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg303_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg856_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg856_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg410_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg656_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg665_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg139_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg142_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg290_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg410_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg118_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg646_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg861_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg421_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg410_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg3_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg687_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg17_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg15_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg11_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg12_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg16_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg8_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg290_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg509_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg789_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg5_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg179_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg15_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg7_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg787_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg403_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg792_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg416_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg508_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg949_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg654_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg533_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg139_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => Delay43No4_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg288_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg503_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg783_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg801_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg416_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg873_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg287_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg546_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg537_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg865_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg664_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg689_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg314_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg326_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg857_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg868_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg424_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add11_3_impl_0_out);

   Delay1No52_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_3_impl_0_out,
                 Y => Delay1No52_out);

SharedReg114_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg114_out;
SharedReg410_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg410_out;
SharedReg143_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg143_out;
SharedReg727_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg727_out;
SharedReg142_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg142_out;
SharedReg141_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg141_out;
SharedReg855_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg855_out;
SharedReg665_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg665_out;
SharedReg931_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg931_out;
SharedReg417_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg417_out;
SharedReg806_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg806_out;
SharedReg805_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg805_out;
SharedReg685_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg685_out;
SharedReg859_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg859_out;
SharedReg285_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg285_out;
SharedReg679_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg679_out;
SharedReg678_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg678_out;
SharedReg803_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg803_out;
SharedReg665_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg665_out;
SharedReg879_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg879_out;
SharedReg160_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg160_out;
SharedReg160_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg160_out;
SharedReg521_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg521_out;
SharedReg139_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg139_out;
SharedReg855_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg855_out;
SharedReg662_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg662_out;
SharedReg519_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg519_out;
SharedReg521_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg521_out;
SharedReg19_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_29_cast <= SharedReg19_out;
SharedReg21_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_30_cast <= SharedReg21_out;
SharedReg35_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_31_cast <= SharedReg35_out;
SharedReg33_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_32_cast <= SharedReg33_out;
SharedReg29_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_33_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_34_cast <= SharedReg30_out;
SharedReg34_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_35_cast <= SharedReg34_out;
SharedReg26_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_36_cast <= SharedReg26_out;
SharedReg289_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_37_cast <= SharedReg289_out;
SharedReg791_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_38_cast <= SharedReg791_out;
SharedReg788_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_39_cast <= SharedReg788_out;
SharedReg23_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_40_cast <= SharedReg23_out;
SharedReg33_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_41_cast <= SharedReg33_out;
SharedReg25_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_42_cast <= SharedReg25_out;
SharedReg503_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_43_cast <= SharedReg503_out;
SharedReg800_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_44_cast <= SharedReg800_out;
SharedReg512_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_45_cast <= SharedReg512_out;
SharedReg526_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_46_cast <= SharedReg526_out;
SharedReg783_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_47_cast <= SharedReg783_out;
SharedReg933_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_48_cast <= SharedReg933_out;
SharedReg676_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_49_cast <= SharedReg676_out;
SharedReg814_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_50_cast <= SharedReg814_out;
SharedReg530_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_51_cast <= SharedReg530_out;
SharedReg283_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_52_cast <= SharedReg283_out;
SharedReg783_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_53_cast <= SharedReg783_out;
SharedReg507_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_54_cast <= SharedReg507_out;
SharedReg526_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_55_cast <= SharedReg526_out;
SharedReg519_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_56_cast <= SharedReg519_out;
SharedReg642_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_57_cast <= SharedReg642_out;
SharedReg161_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_58_cast <= SharedReg161_out;
SharedReg438_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_59_cast <= SharedReg438_out;
SharedReg819_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_60_cast <= SharedReg819_out;
SharedReg684_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_61_cast <= SharedReg684_out;
SharedReg706_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_62_cast <= SharedReg706_out;
SharedReg331_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_63_cast <= SharedReg331_out;
SharedReg285_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_64_cast <= SharedReg285_out;
   MUX_Add11_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg114_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg410_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg806_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg805_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg685_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg859_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg285_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg679_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg678_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg803_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg665_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg879_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg143_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg160_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg160_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg521_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg139_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg855_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg662_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg519_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg521_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg19_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg21_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg727_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg35_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg33_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg29_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg30_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg34_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg26_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg289_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg791_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg788_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg23_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg142_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg33_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg25_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg503_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg800_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg512_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg526_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg783_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg933_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg676_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg814_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg141_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg530_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg283_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg783_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg507_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg526_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg519_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg642_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg161_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg438_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg819_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg855_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg684_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg706_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg331_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg285_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg665_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg931_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg417_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add11_3_impl_1_out);

   Delay1No53_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_3_impl_1_out,
                 Y => Delay1No53_out);

Delay1No54_out_to_Add11_4_impl_parent_implementedSystem_port_0_cast <= Delay1No54_out;
Delay1No55_out_to_Add11_4_impl_parent_implementedSystem_port_1_cast <= Delay1No55_out;
   Add11_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_4_impl_out,
                 X => Delay1No54_out_to_Add11_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No55_out_to_Add11_4_impl_parent_implementedSystem_port_1_cast);

SharedReg431_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg431_out;
SharedReg699_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg699_out;
SharedReg141_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg141_out;
SharedReg997_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg997_out;
SharedReg562_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg562_out;
SharedReg688_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg688_out;
SharedReg711_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg711_out;
SharedReg167_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg167_out;
SharedReg440_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg440_out;
SharedReg142_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg142_out;
SharedReg433_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg433_out;
SharedReg163_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg163_out;
SharedReg985_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg985_out;
SharedReg884_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg884_out;
SharedReg163_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg163_out;
SharedReg695_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg695_out;
SharedReg687_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg687_out;
SharedReg674_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg674_out;
SharedReg439_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg439_out;
SharedReg541_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg541_out;
SharedReg539_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg539_out;
SharedReg882_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg882_out;
SharedReg994_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg994_out;
SharedReg325_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg325_out;
SharedReg686_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg686_out;
SharedReg686_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg686_out;
SharedReg425_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg425_out;
SharedReg432_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg432_out;
SharedReg711_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_29_cast <= SharedReg711_out;
SharedReg168_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_30_cast <= SharedReg168_out;
SharedReg315_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_31_cast <= SharedReg315_out;
SharedReg425_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_32_cast <= SharedReg425_out;
SharedReg142_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_33_cast <= SharedReg142_out;
SharedReg667_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_34_cast <= SharedReg667_out;
SharedReg691_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_35_cast <= SharedReg691_out;
SharedReg436_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_36_cast <= SharedReg436_out;
SharedReg425_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_37_cast <= SharedReg425_out;
SharedReg1_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1_out;
SharedReg3_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_39_cast <= SharedReg3_out;
SharedReg172_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_40_cast <= SharedReg172_out;
SharedReg191_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_41_cast <= SharedReg191_out;
SharedReg824_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_42_cast <= SharedReg824_out;
SharedReg12_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_43_cast <= SharedReg12_out;
SharedReg16_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_44_cast <= SharedReg16_out;
SharedReg8_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_45_cast <= SharedReg8_out;
SharedReg315_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_46_cast <= SharedReg315_out;
SharedReg525_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_47_cast <= SharedReg525_out;
SharedReg807_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_48_cast <= SharedReg807_out;
SharedReg5_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_49_cast <= SharedReg5_out;
SharedReg15_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_50_cast <= SharedReg15_out;
SharedReg11_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_51_cast <= SharedReg11_out;
SharedReg805_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_52_cast <= SharedReg805_out;
SharedReg418_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_53_cast <= SharedReg418_out;
SharedReg810_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_54_cast <= SharedReg810_out;
SharedReg827_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_55_cast <= SharedReg827_out;
SharedReg431_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_56_cast <= SharedReg431_out;
SharedReg172_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_57_cast <= SharedReg172_out;
SharedReg716_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_58_cast <= SharedReg716_out;
SharedReg5_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_59_cast <= SharedReg5_out;
SharedReg4_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_60_cast <= SharedReg4_out;
SharedReg836_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_61_cast <= SharedReg836_out;
SharedReg425_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_62_cast <= SharedReg425_out;
SharedReg425_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_63_cast <= SharedReg425_out;
SharedReg13_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_64_cast <= SharedReg13_out;
   MUX_Add11_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg431_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg699_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg433_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg163_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg985_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg884_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg163_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg695_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg687_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg674_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg439_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg541_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg141_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg539_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg882_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg994_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg325_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg686_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg686_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg425_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg432_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg711_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg168_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg997_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg315_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg425_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg142_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg667_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg691_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg436_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg425_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg3_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg172_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg562_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg191_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg824_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg12_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg16_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg8_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg315_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg525_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg807_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg5_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg15_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg688_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg11_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg805_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg418_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg810_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg827_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg431_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg172_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg716_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg5_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg4_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg711_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg836_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg425_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg425_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg13_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg167_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg440_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg142_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add11_4_impl_0_out);

   Delay1No54_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_4_impl_0_out,
                 Y => Delay1No54_out);

SharedReg535_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg535_out;
SharedReg857_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg857_out;
SharedReg330_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg330_out;
SharedReg996_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg996_out;
SharedReg453_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg453_out;
SharedReg705_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg705_out;
SharedReg728_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg728_out;
SharedReg185_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg185_out;
SharedReg447_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg447_out;
SharedReg139_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg139_out;
SharedReg425_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg425_out;
SharedReg169_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg169_out;
SharedReg904_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg904_out;
SharedReg1001_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1001_out;
SharedReg165_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg165_out;
SharedReg685_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg685_out;
SharedReg711_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg711_out;
SharedReg855_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg855_out;
SharedReg432_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg432_out;
SharedReg824_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg824_out;
SharedReg823_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg823_out;
SharedReg712_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg712_out;
SharedReg685_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg685_out;
SharedReg310_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg310_out;
SharedReg723_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg723_out;
SharedReg722_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg722_out;
SharedReg821_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg821_out;
SharedReg425_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg425_out;
SharedReg702_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_29_cast <= SharedReg702_out;
SharedReg183_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_30_cast <= SharedReg183_out;
SharedReg183_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_31_cast <= SharedReg183_out;
SharedReg537_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_32_cast <= SharedReg537_out;
SharedReg310_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_33_cast <= SharedReg310_out;
SharedReg685_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_34_cast <= SharedReg685_out;
SharedReg708_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_35_cast <= SharedReg708_out;
SharedReg535_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_36_cast <= SharedReg535_out;
SharedReg537_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_37_cast <= SharedReg537_out;
SharedReg19_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_38_cast <= SharedReg19_out;
SharedReg21_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_39_cast <= SharedReg21_out;
SharedReg163_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_40_cast <= SharedReg163_out;
SharedReg348_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_41_cast <= SharedReg348_out;
SharedReg826_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_42_cast <= SharedReg826_out;
SharedReg30_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_43_cast <= SharedReg30_out;
SharedReg34_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_44_cast <= SharedReg34_out;
SharedReg26_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_45_cast <= SharedReg26_out;
SharedReg314_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_46_cast <= SharedReg314_out;
SharedReg809_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_47_cast <= SharedReg809_out;
SharedReg806_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_48_cast <= SharedReg806_out;
SharedReg23_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_49_cast <= SharedReg23_out;
SharedReg33_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_50_cast <= SharedReg33_out;
SharedReg29_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_51_cast <= SharedReg29_out;
SharedReg519_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_52_cast <= SharedReg519_out;
SharedReg818_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_53_cast <= SharedReg818_out;
SharedReg528_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_54_cast <= SharedReg528_out;
SharedReg543_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_55_cast <= SharedReg543_out;
SharedReg539_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_56_cast <= SharedReg539_out;
SharedReg318_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_57_cast <= SharedReg318_out;
SharedReg696_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_58_cast <= SharedReg696_out;
SharedReg23_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_59_cast <= SharedReg23_out;
SharedReg22_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_60_cast <= SharedReg22_out;
SharedReg434_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_61_cast <= SharedReg434_out;
SharedReg535_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_62_cast <= SharedReg535_out;
SharedReg432_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_63_cast <= SharedReg432_out;
SharedReg31_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_64_cast <= SharedReg31_out;
   MUX_Add11_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg535_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg857_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg425_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg169_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg904_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1001_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg165_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg685_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg711_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg855_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg432_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg824_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg330_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg823_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg712_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg685_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg310_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg723_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg722_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg821_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg425_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg702_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg183_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg996_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg183_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg537_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg310_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg685_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg708_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg535_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg537_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg19_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg21_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg163_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg453_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg348_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg826_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg30_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg34_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg26_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg314_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg809_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg806_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg23_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg33_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg705_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg29_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg519_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg818_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg528_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg543_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg539_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg318_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg696_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg23_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg22_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg728_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg434_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg535_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg432_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg31_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg185_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg447_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg139_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Add11_4_impl_1_out);

   Delay1No55_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_4_impl_1_out,
                 Y => Delay1No55_out);

Delay1No56_out_to_Add11_6_impl_parent_implementedSystem_port_0_cast <= Delay1No56_out;
Delay1No57_out_to_Add11_6_impl_parent_implementedSystem_port_1_cast <= Delay1No57_out;
   Add11_6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_6_impl_out,
                 X => Delay1No56_out_to_Add11_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No57_out_to_Add11_6_impl_parent_implementedSystem_port_1_cast);

SharedReg1_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1_out;
SharedReg11_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg11_out;
SharedReg12_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg12_out;
SharedReg16_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg16_out;
SharedReg717_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg717_out;
SharedReg199_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg199_out;
SharedReg551_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg551_out;
SharedReg440_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg440_out;
SharedReg556_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg556_out;
SharedReg454_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg454_out;
SharedReg440_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg440_out;
SharedReg447_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg447_out;
SharedReg337_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_13_cast <= SharedReg337_out;
SharedReg440_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_14_cast <= SharedReg440_out;
SharedReg844_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_15_cast <= SharedReg844_out;
SharedReg888_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_16_cast <= SharedReg888_out;
SharedReg335_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_17_cast <= SharedReg335_out;
SharedReg843_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_18_cast <= SharedReg843_out;
SharedReg440_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_19_cast <= SharedReg440_out;
SharedReg842_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_20_cast <= SharedReg842_out;
SharedReg551_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_21_cast <= SharedReg551_out;
Delay43No6_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_22_cast <= Delay43No6_out;
SharedReg448_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_23_cast <= SharedReg448_out;
SharedReg557_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_24_cast <= SharedReg557_out;
SharedReg333_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_25_cast <= SharedReg333_out;
SharedReg566_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_26_cast <= SharedReg566_out;
SharedReg442_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_27_cast <= SharedReg442_out;
SharedReg845_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_28_cast <= SharedReg845_out;
SharedReg446_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_29_cast <= SharedReg446_out;
SharedReg839_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_30_cast <= SharedReg839_out;
SharedReg342_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_31_cast <= SharedReg342_out;
SharedReg841_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_32_cast <= SharedReg841_out;
SharedReg837_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_33_cast <= SharedReg837_out;
   MUX_Add11_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_33_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg11_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg440_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg447_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg337_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg440_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg844_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg888_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg335_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg843_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg440_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg842_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg12_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg551_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => Delay43No6_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg448_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg557_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg333_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg566_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg442_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg845_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg446_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg839_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg16_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg342_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg841_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg837_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_33_cast,
                 iS_4 => SharedReg717_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg199_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg551_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg440_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg556_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg454_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Add11_6_impl_0_LUT_out,
                 oMux => MUX_Add11_6_impl_0_out);

   Delay1No56_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_6_impl_0_out,
                 Y => Delay1No56_out);

SharedReg19_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg19_out;
SharedReg29_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg30_out;
SharedReg34_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg34_out;
SharedReg837_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg837_out;
SharedReg552_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg552_out;
SharedReg186_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg186_out;
SharedReg837_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg837_out;
SharedReg553_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg553_out;
SharedReg440_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg440_out;
SharedReg555_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg555_out;
SharedReg839_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg839_out;
SharedReg441_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_13_cast <= SharedReg441_out;
SharedReg837_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_14_cast <= SharedReg837_out;
SharedReg882_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_15_cast <= SharedReg882_out;
SharedReg841_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_16_cast <= SharedReg841_out;
SharedReg844_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_17_cast <= SharedReg844_out;
SharedReg332_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_18_cast <= SharedReg332_out;
SharedReg845_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_19_cast <= SharedReg845_out;
SharedReg562_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_20_cast <= SharedReg562_out;
SharedReg854_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_21_cast <= SharedReg854_out;
SharedReg207_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_22_cast <= SharedReg207_out;
SharedReg845_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_23_cast <= SharedReg845_out;
SharedReg842_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_24_cast <= SharedReg842_out;
SharedReg346_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_25_cast <= SharedReg346_out;
SharedReg551_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_26_cast <= SharedReg551_out;
SharedReg983_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_27_cast <= SharedReg983_out;
SharedReg559_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_28_cast <= SharedReg559_out;
SharedReg444_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_29_cast <= SharedReg444_out;
SharedReg838_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_30_cast <= SharedReg838_out;
SharedReg186_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_31_cast <= SharedReg186_out;
SharedReg558_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_32_cast <= SharedReg558_out;
SharedReg551_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_33_cast <= SharedReg551_out;
   MUX_Add11_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_33_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg19_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg29_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg555_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg839_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg441_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg837_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg882_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg841_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg844_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg332_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg845_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg562_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg30_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg854_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg207_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg845_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg842_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg346_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg551_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg983_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg559_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg444_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg838_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg34_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg186_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg558_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg551_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_33_cast,
                 iS_4 => SharedReg837_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg552_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg186_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg837_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg553_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg440_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Add11_6_impl_1_LUT_out,
                 oMux => MUX_Add11_6_impl_1_out);

   Delay1No57_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_6_impl_1_out,
                 Y => Delay1No57_out);

Delay1No58_out_to_Product4_0_impl_parent_implementedSystem_port_0_cast <= Delay1No58_out;
Delay1No59_out_to_Product4_0_impl_parent_implementedSystem_port_1_cast <= Delay1No59_out;
   Product4_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_0_impl_out,
                 X => Delay1No58_out_to_Product4_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No59_out_to_Product4_0_impl_parent_implementedSystem_port_1_cast);

SharedReg1044_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1044_out;
SharedReg1045_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1045_out;
SharedReg1104_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1104_out;
SharedReg1055_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1055_out;
SharedReg1056_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1056_out;
SharedReg977_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg977_out;
SharedReg1057_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1057_out;
SharedReg1003_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1003_out;
SharedReg957_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg957_out;
SharedReg1108_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1108_out;
SharedReg1154_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1154_out;
SharedReg570_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg570_out;
SharedReg1007_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1007_out;
SharedReg1008_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1008_out;
SharedReg962_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg962_out;
SharedReg1010_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1010_out;
SharedReg1150_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1150_out;
SharedReg1011_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1011_out;
SharedReg1123_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1123_out;
SharedReg1124_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1124_out;
SharedReg574_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg574_out;
SharedReg1120_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1120_out;
SharedReg968_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg968_out;
SharedReg1151_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1151_out;
SharedReg1016_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1016_out;
SharedReg1068_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1068_out;
SharedReg1161_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1161_out;
SharedReg1155_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1155_out;
SharedReg1048_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1048_out;
SharedReg1049_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1049_out;
SharedReg1099_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1099_out;
SharedReg1051_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1051_out;
SharedReg1052_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1052_out;
SharedReg1019_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1019_out;
SharedReg1020_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1020_out;
SharedReg1021_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1021_out;
SharedReg1022_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1022_out;
SharedReg1023_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1023_out;
SharedReg1111_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1111_out;
SharedReg1024_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1024_out;
SharedReg1025_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1025_out;
SharedReg1113_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1113_out;
SharedReg1076_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1076_out;
SharedReg1027_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1027_out;
SharedReg1028_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1028_out;
SharedReg1029_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1029_out;
SharedReg1030_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1030_out;
SharedReg1031_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1031_out;
SharedReg1080_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1080_out;
SharedReg1032_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1032_out;
SharedReg1033_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1033_out;
SharedReg1034_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1034_out;
SharedReg1035_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1035_out;
SharedReg1085_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1085_out;
SharedReg49_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_55_cast <= SharedReg49_out;
SharedReg1054_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1054_out;
SharedReg1038_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1038_out;
SharedReg1039_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1039_out;
SharedReg1040_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1040_out;
SharedReg1041_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1041_out;
SharedReg1130_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1130_out;
SharedReg1042_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1042_out;
SharedReg36_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_63_cast <= SharedReg36_out;
SharedReg1043_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1043_out;
   MUX_Product4_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1044_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1045_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1154_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg570_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1007_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1008_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg962_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1010_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1150_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1011_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1123_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1124_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1104_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg574_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1120_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg968_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1151_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1016_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1068_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1161_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1155_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1048_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1049_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1055_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1099_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1051_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1052_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1019_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1020_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1021_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1022_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1023_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1111_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1024_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1056_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1025_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1113_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1076_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1027_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1028_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1029_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1030_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1031_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1080_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1032_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg977_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1033_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1034_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1035_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1085_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg49_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1054_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1038_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1039_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1040_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1041_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1057_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1130_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1042_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg36_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1043_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1003_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg957_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1108_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product4_0_impl_0_out);

   Delay1No58_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_0_impl_0_out,
                 Y => Delay1No58_out);

SharedReg37_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg37_out;
SharedReg37_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg37_out;
SharedReg978_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg978_out;
SharedReg980_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg980_out;
SharedReg57_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg57_out;
SharedReg1107_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1107_out;
SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg36_out;
SharedReg37_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg37_out;
SharedReg1168_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1168_out;
SharedReg957_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg957_out;
SharedReg569_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg569_out;
SharedReg1160_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1160_out;
SharedReg213_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg213_out;
SharedReg215_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg215_out;
SharedReg1114_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1114_out;
SharedReg44_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg44_out;
SharedReg963_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg963_out;
SharedReg42_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg42_out;
SharedReg573_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg573_out;
SharedReg575_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg575_out;
SharedReg1121_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1121_out;
SharedReg577_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg577_out;
SharedReg1153_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1153_out;
SharedReg969_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg969_out;
SharedReg219_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg219_out;
SharedReg49_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg49_out;
SharedReg970_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg970_out;
SharedReg971_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg971_out;
SharedReg48_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_29_cast <= SharedReg48_out;
SharedReg48_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_30_cast <= SharedReg48_out;
SharedReg221_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_31_cast <= SharedReg221_out;
SharedReg222_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_32_cast <= SharedReg222_out;
SharedReg45_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_33_cast <= SharedReg45_out;
SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_34_cast <= SharedReg36_out;
SharedReg957_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_35_cast <= SharedReg957_out;
SharedReg208_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_36_cast <= SharedReg208_out;
SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_37_cast <= SharedReg36_out;
SharedReg208_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_38_cast <= SharedReg208_out;
SharedReg958_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_39_cast <= SharedReg958_out;
SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_40_cast <= SharedReg36_out;
SharedReg209_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_41_cast <= SharedReg209_out;
SharedReg958_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_42_cast <= SharedReg958_out;
SharedReg43_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_43_cast <= SharedReg43_out;
SharedReg44_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_44_cast <= SharedReg44_out;
SharedReg214_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_45_cast <= SharedReg214_out;
SharedReg964_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_46_cast <= SharedReg964_out;
SharedReg214_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_47_cast <= SharedReg214_out;
SharedReg43_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_48_cast <= SharedReg43_out;
SharedReg44_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_49_cast <= SharedReg44_out;
SharedReg216_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_50_cast <= SharedReg216_out;
SharedReg49_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_51_cast <= SharedReg49_out;
SharedReg40_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_52_cast <= SharedReg40_out;
SharedReg580_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_53_cast <= SharedReg580_out;
SharedReg38_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_54_cast <= SharedReg38_out;
SharedReg1086_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_55_cast <= SharedReg1086_out;
SharedReg56_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_56_cast <= SharedReg56_out;
SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_57_cast <= SharedReg36_out;
SharedReg208_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_58_cast <= SharedReg208_out;
SharedReg37_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_59_cast <= SharedReg37_out;
SharedReg37_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_60_cast <= SharedReg37_out;
SharedReg570_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_61_cast <= SharedReg570_out;
SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_62_cast <= SharedReg36_out;
SharedReg1092_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_63_cast <= SharedReg1092_out;
SharedReg37_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_64_cast <= SharedReg37_out;
   MUX_Product4_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg37_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg37_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg569_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1160_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg213_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg215_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1114_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg44_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg963_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg42_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg573_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg575_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg978_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1121_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg577_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1153_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg969_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg219_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg49_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg970_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg971_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg48_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg48_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg980_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg221_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg222_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg45_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg957_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg208_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg208_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg958_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg57_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg209_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg958_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg43_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg44_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg214_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg964_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg214_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg43_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg44_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg216_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1107_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg49_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg40_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg580_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg38_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1086_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg56_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg208_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg37_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg37_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg570_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1092_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg37_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg37_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1168_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg957_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product4_0_impl_1_out);

   Delay1No59_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_0_impl_1_out,
                 Y => Delay1No59_out);

Delay1No60_out_to_Product4_1_impl_parent_implementedSystem_port_0_cast <= Delay1No60_out;
Delay1No61_out_to_Product4_1_impl_parent_implementedSystem_port_1_cast <= Delay1No61_out;
   Product4_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_1_impl_out,
                 X => Delay1No60_out_to_Product4_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No61_out_to_Product4_1_impl_parent_implementedSystem_port_1_cast);

SharedReg1054_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1054_out;
SharedReg1038_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1038_out;
SharedReg1039_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1039_out;
SharedReg1040_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1040_out;
SharedReg1041_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1041_out;
SharedReg1130_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1130_out;
SharedReg1042_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1042_out;
SharedReg62_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg62_out;
SharedReg1043_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1043_out;
SharedReg1044_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1044_out;
SharedReg1045_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1045_out;
SharedReg1104_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1104_out;
SharedReg1055_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1055_out;
SharedReg1056_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1056_out;
SharedReg925_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg925_out;
SharedReg1057_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1057_out;
SharedReg1003_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1003_out;
SharedReg906_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg906_out;
SharedReg1108_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1108_out;
SharedReg1154_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1154_out;
SharedReg596_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg596_out;
SharedReg1007_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1007_out;
SharedReg1008_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1008_out;
SharedReg911_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg911_out;
SharedReg1010_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1010_out;
SharedReg1150_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1150_out;
SharedReg1011_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1011_out;
SharedReg1123_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1123_out;
SharedReg1124_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1124_out;
SharedReg964_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_30_cast <= SharedReg964_out;
SharedReg1120_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1120_out;
SharedReg917_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_32_cast <= SharedReg917_out;
SharedReg1151_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1151_out;
SharedReg1016_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1016_out;
SharedReg1068_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1068_out;
SharedReg1161_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1161_out;
SharedReg1155_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1155_out;
SharedReg1048_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1048_out;
SharedReg1049_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1049_out;
SharedReg1099_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1099_out;
SharedReg1051_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1051_out;
SharedReg1052_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1052_out;
SharedReg1019_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1019_out;
SharedReg1020_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1020_out;
SharedReg1021_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1021_out;
SharedReg1022_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1022_out;
SharedReg1023_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1023_out;
SharedReg1111_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1111_out;
SharedReg1024_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1024_out;
SharedReg1025_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1025_out;
SharedReg1113_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1113_out;
SharedReg1076_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1076_out;
SharedReg1027_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1027_out;
SharedReg1028_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1028_out;
SharedReg1029_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1029_out;
SharedReg1030_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1030_out;
SharedReg1031_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1031_out;
SharedReg1080_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1080_out;
SharedReg1032_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1032_out;
SharedReg1033_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1033_out;
SharedReg1034_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1034_out;
SharedReg1035_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1035_out;
SharedReg1085_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1085_out;
SharedReg75_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_64_cast <= SharedReg75_out;
   MUX_Product4_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1054_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1038_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1045_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1104_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1055_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1056_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg925_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1057_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1003_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg906_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1108_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1154_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1039_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg596_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1007_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1008_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg911_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1010_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1150_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1011_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1123_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1124_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg964_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1040_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1120_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg917_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1151_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1016_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1068_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1161_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1155_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1048_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1049_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1099_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1041_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1051_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1052_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1019_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1020_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1021_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1022_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1023_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1111_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1024_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1025_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1130_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1113_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1076_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1027_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1028_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1029_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1030_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1031_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1080_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1032_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1033_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1042_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1034_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1035_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1085_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg75_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg62_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1043_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1044_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product4_1_impl_0_out);

   Delay1No60_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_1_impl_0_out,
                 Y => Delay1No60_out);

SharedReg80_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg80_out;
SharedReg208_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg208_out;
SharedReg62_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg62_out;
SharedReg209_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg209_out;
SharedReg209_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg209_out;
SharedReg960_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg960_out;
SharedReg62_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg62_out;
SharedReg1092_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1092_out;
SharedReg63_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg63_out;
SharedReg63_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg63_out;
SharedReg63_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg63_out;
SharedReg926_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg926_out;
SharedReg928_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg928_out;
SharedReg83_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg83_out;
SharedReg1107_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1107_out;
SharedReg62_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg62_out;
SharedReg63_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg63_out;
SharedReg1168_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1168_out;
SharedReg906_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg906_out;
SharedReg595_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg595_out;
SharedReg1160_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1160_out;
SharedReg239_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg239_out;
SharedReg241_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg241_out;
SharedReg1114_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1114_out;
SharedReg70_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg70_out;
SharedReg912_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg912_out;
SharedReg68_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg68_out;
SharedReg599_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg599_out;
SharedReg601_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_29_cast <= SharedReg601_out;
SharedReg1121_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_30_cast <= SharedReg1121_out;
SharedReg603_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_31_cast <= SharedReg603_out;
SharedReg1153_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_32_cast <= SharedReg1153_out;
SharedReg918_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_33_cast <= SharedReg918_out;
SharedReg245_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_34_cast <= SharedReg245_out;
SharedReg75_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_35_cast <= SharedReg75_out;
SharedReg605_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_36_cast <= SharedReg605_out;
SharedReg606_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_37_cast <= SharedReg606_out;
SharedReg74_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_38_cast <= SharedReg74_out;
SharedReg74_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_39_cast <= SharedReg74_out;
SharedReg247_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_40_cast <= SharedReg247_out;
SharedReg248_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_41_cast <= SharedReg248_out;
SharedReg217_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_42_cast <= SharedReg217_out;
SharedReg62_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_43_cast <= SharedReg62_out;
SharedReg906_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_44_cast <= SharedReg906_out;
SharedReg62_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_45_cast <= SharedReg62_out;
SharedReg36_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_46_cast <= SharedReg36_out;
SharedReg62_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_47_cast <= SharedReg62_out;
SharedReg594_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_48_cast <= SharedReg594_out;
SharedReg62_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_49_cast <= SharedReg62_out;
SharedReg235_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_50_cast <= SharedReg235_out;
SharedReg907_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_51_cast <= SharedReg907_out;
SharedReg215_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_52_cast <= SharedReg215_out;
SharedReg216_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_53_cast <= SharedReg216_out;
SharedReg240_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_54_cast <= SharedReg240_out;
SharedReg913_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_55_cast <= SharedReg913_out;
SharedReg240_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_56_cast <= SharedReg240_out;
SharedReg69_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_57_cast <= SharedReg69_out;
SharedReg70_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_58_cast <= SharedReg70_out;
SharedReg242_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_59_cast <= SharedReg242_out;
SharedReg221_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_60_cast <= SharedReg221_out;
SharedReg66_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_61_cast <= SharedReg66_out;
SharedReg972_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_62_cast <= SharedReg972_out;
SharedReg210_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_63_cast <= SharedReg210_out;
SharedReg1086_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_64_cast <= SharedReg1086_out;
   MUX_Product4_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg80_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg208_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg63_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg926_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg928_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg83_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1107_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg62_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg63_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1168_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg906_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg595_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg62_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1160_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg239_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg241_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1114_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg70_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg912_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg68_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg599_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg601_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1121_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg209_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg603_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1153_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg918_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg245_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg75_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg605_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg606_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg74_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg74_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg247_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg209_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg248_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg217_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg62_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg906_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg62_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg36_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg62_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg594_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg62_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg235_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg960_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg907_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg215_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg216_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg240_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg913_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg240_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg69_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg70_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg242_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg221_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg62_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg66_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg972_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg210_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1086_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1092_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg63_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg63_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product4_1_impl_1_out);

   Delay1No61_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_1_impl_1_out,
                 Y => Delay1No61_out);

Delay1No62_out_to_Product4_2_impl_parent_implementedSystem_port_0_cast <= Delay1No62_out;
Delay1No63_out_to_Product4_2_impl_parent_implementedSystem_port_1_cast <= Delay1No63_out;
   Product4_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_2_impl_out,
                 X => Delay1No62_out_to_Product4_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No63_out_to_Product4_2_impl_parent_implementedSystem_port_1_cast);

SharedReg1030_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1030_out;
SharedReg1031_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1031_out;
SharedReg1080_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1080_out;
SharedReg1032_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1032_out;
SharedReg1033_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1033_out;
SharedReg1034_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1034_out;
SharedReg1035_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1035_out;
SharedReg1085_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1085_out;
SharedReg247_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg247_out;
SharedReg1054_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1054_out;
SharedReg1038_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1038_out;
SharedReg1039_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1039_out;
SharedReg1040_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1040_out;
SharedReg1041_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1041_out;
SharedReg1130_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1130_out;
SharedReg1042_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1042_out;
SharedReg88_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg88_out;
SharedReg1043_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1043_out;
SharedReg1044_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1044_out;
SharedReg1045_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1045_out;
SharedReg1104_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1104_out;
SharedReg1055_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1055_out;
SharedReg1056_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1056_out;
SharedReg951_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg951_out;
SharedReg1057_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1057_out;
SharedReg1003_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1003_out;
SharedReg931_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg931_out;
SharedReg1108_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1108_out;
SharedReg1154_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1154_out;
SharedReg620_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_30_cast <= SharedReg620_out;
SharedReg1007_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1007_out;
SharedReg1008_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1008_out;
SharedReg936_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_33_cast <= SharedReg936_out;
SharedReg1010_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1010_out;
SharedReg1150_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1150_out;
SharedReg1011_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1011_out;
SharedReg1123_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1123_out;
SharedReg1124_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1124_out;
SharedReg913_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_39_cast <= SharedReg913_out;
SharedReg1120_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1120_out;
SharedReg942_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_41_cast <= SharedReg942_out;
SharedReg1151_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1151_out;
SharedReg1016_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1016_out;
SharedReg1068_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1068_out;
SharedReg1161_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1161_out;
SharedReg1155_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1155_out;
SharedReg1048_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1048_out;
SharedReg1049_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1049_out;
SharedReg1099_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1099_out;
SharedReg1051_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1051_out;
SharedReg1052_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1052_out;
SharedReg1019_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1019_out;
SharedReg1020_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1020_out;
SharedReg1021_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1021_out;
SharedReg1022_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1022_out;
SharedReg1023_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1023_out;
SharedReg1111_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1111_out;
SharedReg1024_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1024_out;
SharedReg1025_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1025_out;
SharedReg1113_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1113_out;
SharedReg1076_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1076_out;
SharedReg1027_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1027_out;
SharedReg1028_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1028_out;
SharedReg1029_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1029_out;
   MUX_Product4_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1030_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1031_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1038_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1039_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1040_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1041_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1130_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1042_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg88_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1043_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1044_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1045_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1080_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1104_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1055_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1056_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg951_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1057_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1003_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg931_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1108_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1154_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg620_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1032_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1007_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1008_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg936_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1010_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1150_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1011_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1123_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1124_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg913_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1120_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1033_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg942_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1151_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1016_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1068_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1161_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1155_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1048_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1049_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1099_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1051_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1034_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1052_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1019_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1020_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1021_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1022_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1023_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1111_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1024_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1025_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1113_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1035_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1076_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1027_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1028_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1029_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1085_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg247_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1054_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product4_2_impl_0_out);

   Delay1No62_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_2_impl_0_out,
                 Y => Delay1No62_out);

SharedReg266_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg266_out;
SharedReg94_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg94_out;
SharedReg95_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg95_out;
SharedReg95_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg95_out;
SharedReg75_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg75_out;
SharedReg238_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg238_out;
SharedReg607_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg607_out;
SharedReg236_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg236_out;
SharedReg1086_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1086_out;
SharedReg105_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg105_out;
SharedReg234_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg234_out;
SharedReg88_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg88_out;
SharedReg235_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg235_out;
SharedReg235_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg235_out;
SharedReg909_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg909_out;
SharedReg88_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg88_out;
SharedReg1092_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1092_out;
SharedReg89_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg89_out;
SharedReg89_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg89_out;
SharedReg89_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg89_out;
SharedReg952_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg952_out;
SharedReg954_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg954_out;
SharedReg255_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg255_out;
SharedReg1107_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1107_out;
SharedReg88_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg88_out;
SharedReg89_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg89_out;
SharedReg1168_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1168_out;
SharedReg931_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg931_out;
SharedReg619_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_29_cast <= SharedReg619_out;
SharedReg1160_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_30_cast <= SharedReg1160_out;
SharedReg265_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_31_cast <= SharedReg265_out;
SharedReg267_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_32_cast <= SharedReg267_out;
SharedReg1114_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_33_cast <= SharedReg1114_out;
SharedReg95_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_34_cast <= SharedReg95_out;
SharedReg937_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_35_cast <= SharedReg937_out;
SharedReg93_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_36_cast <= SharedReg93_out;
SharedReg623_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_37_cast <= SharedReg623_out;
SharedReg625_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_38_cast <= SharedReg625_out;
SharedReg1121_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_39_cast <= SharedReg1121_out;
SharedReg628_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_40_cast <= SharedReg628_out;
SharedReg1153_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_41_cast <= SharedReg1153_out;
SharedReg943_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_42_cast <= SharedReg943_out;
SharedReg271_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_43_cast <= SharedReg271_out;
SharedReg100_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_44_cast <= SharedReg100_out;
SharedReg630_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_45_cast <= SharedReg630_out;
SharedReg631_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_46_cast <= SharedReg631_out;
SharedReg99_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_47_cast <= SharedReg99_out;
SharedReg99_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_48_cast <= SharedReg99_out;
SharedReg273_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_49_cast <= SharedReg273_out;
SharedReg274_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_50_cast <= SharedReg274_out;
SharedReg243_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_51_cast <= SharedReg243_out;
SharedReg88_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_52_cast <= SharedReg88_out;
SharedReg931_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_53_cast <= SharedReg931_out;
SharedReg88_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_54_cast <= SharedReg88_out;
SharedReg62_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_55_cast <= SharedReg62_out;
SharedReg234_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_56_cast <= SharedReg234_out;
SharedReg907_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_57_cast <= SharedReg907_out;
SharedReg88_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_58_cast <= SharedReg88_out;
SharedReg261_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_59_cast <= SharedReg261_out;
SharedReg932_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_60_cast <= SharedReg932_out;
SharedReg241_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_61_cast <= SharedReg241_out;
SharedReg242_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_62_cast <= SharedReg242_out;
SharedReg266_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_63_cast <= SharedReg266_out;
SharedReg938_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_64_cast <= SharedReg938_out;
   MUX_Product4_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg266_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg94_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg234_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg88_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg235_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg235_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg909_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg88_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1092_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg89_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg89_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg89_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg95_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg952_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg954_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg255_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1107_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg88_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg89_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1168_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg931_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg619_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1160_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg95_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg265_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg267_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1114_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg95_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg937_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg93_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg623_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg625_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1121_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg628_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg75_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1153_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg943_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg271_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg100_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg630_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg631_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg99_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg99_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg273_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg274_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg238_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg243_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg88_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg931_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg88_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg62_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg234_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg907_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg88_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg261_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg932_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg607_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg241_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg242_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg266_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg938_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg236_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1086_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg105_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product4_2_impl_1_out);

   Delay1No63_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_2_impl_1_out,
                 Y => Delay1No63_out);

Delay1No64_out_to_Product4_3_impl_parent_implementedSystem_port_0_cast <= Delay1No64_out;
Delay1No65_out_to_Product4_3_impl_parent_implementedSystem_port_1_cast <= Delay1No65_out;
   Product4_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_3_impl_out,
                 X => Delay1No64_out_to_Product4_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No65_out_to_Product4_3_impl_parent_implementedSystem_port_1_cast);

SharedReg1023_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1023_out;
SharedReg1111_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1111_out;
SharedReg1024_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1024_out;
SharedReg1025_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1025_out;
SharedReg1113_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1113_out;
SharedReg1076_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1076_out;
SharedReg1027_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1027_out;
SharedReg1028_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1028_out;
SharedReg1029_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1029_out;
SharedReg1030_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1030_out;
SharedReg1031_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1031_out;
SharedReg1080_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1080_out;
SharedReg1032_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1032_out;
SharedReg1033_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1033_out;
SharedReg1034_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1034_out;
SharedReg1035_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1035_out;
SharedReg1085_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1085_out;
SharedReg100_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg100_out;
SharedReg1054_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1054_out;
SharedReg1038_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1038_out;
SharedReg1039_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1039_out;
SharedReg1040_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1040_out;
SharedReg1041_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1041_out;
SharedReg1130_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1130_out;
SharedReg1042_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1042_out;
SharedReg114_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg114_out;
SharedReg1043_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1043_out;
SharedReg1044_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1044_out;
SharedReg1045_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1045_out;
SharedReg1104_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1104_out;
SharedReg1055_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1055_out;
SharedReg1056_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1056_out;
SharedReg876_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_33_cast <= SharedReg876_out;
SharedReg1057_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1057_out;
SharedReg1003_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1003_out;
SharedReg855_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_36_cast <= SharedReg855_out;
SharedReg1108_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1108_out;
SharedReg1154_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1154_out;
SharedReg643_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_39_cast <= SharedReg643_out;
SharedReg1007_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1007_out;
SharedReg1008_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1008_out;
SharedReg860_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_42_cast <= SharedReg860_out;
SharedReg1010_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1010_out;
SharedReg1150_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1150_out;
SharedReg1011_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1011_out;
SharedReg1123_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1123_out;
SharedReg1124_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1124_out;
SharedReg938_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_48_cast <= SharedReg938_out;
SharedReg1120_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1120_out;
SharedReg866_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_50_cast <= SharedReg866_out;
SharedReg1151_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1151_out;
SharedReg1016_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1016_out;
SharedReg1068_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1068_out;
SharedReg1161_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1161_out;
SharedReg1155_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1155_out;
SharedReg1048_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1048_out;
SharedReg1049_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1049_out;
SharedReg1099_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1099_out;
SharedReg1051_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1051_out;
SharedReg1052_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1052_out;
SharedReg1019_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1019_out;
SharedReg1020_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1020_out;
SharedReg1021_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1021_out;
SharedReg1022_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1022_out;
   MUX_Product4_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1023_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1111_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1031_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1080_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1032_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1033_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1034_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1035_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1085_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg100_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1054_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1038_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1024_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1039_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1040_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1041_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1130_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1042_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg114_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1043_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1044_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1045_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1104_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1025_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1055_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1056_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg876_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1057_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1003_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg855_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1108_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1154_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg643_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1007_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1113_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1008_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg860_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1010_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1150_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1011_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1123_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1124_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg938_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1120_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg866_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1076_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1151_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1016_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1068_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1161_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1155_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1048_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1049_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1099_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1051_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1052_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1027_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1019_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1020_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1021_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1022_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1028_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1029_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1030_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product4_3_impl_0_out);

   Delay1No64_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_3_impl_0_out,
                 Y => Delay1No64_out);

SharedReg88_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg88_out;
SharedReg618_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg618_out;
SharedReg260_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg260_out;
SharedReg115_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg115_out;
SharedReg641_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg641_out;
SharedReg94_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg94_out;
SharedReg95_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg95_out;
SharedReg119_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg119_out;
SharedReg647_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg647_out;
SharedReg119_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg119_out;
SharedReg267_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg267_out;
SharedReg268_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg268_out;
SharedReg268_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg268_out;
SharedReg247_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg247_out;
SharedReg264_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg264_out;
SharedReg920_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg920_out;
SharedReg262_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg262_out;
SharedReg1086_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1086_out;
SharedReg130_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg130_out;
SharedReg260_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg260_out;
SharedReg114_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg114_out;
SharedReg261_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg261_out;
SharedReg261_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg261_out;
SharedReg934_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg934_out;
SharedReg114_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg114_out;
SharedReg1092_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1092_out;
SharedReg115_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg115_out;
SharedReg115_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg115_out;
SharedReg115_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_29_cast <= SharedReg115_out;
SharedReg877_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_30_cast <= SharedReg877_out;
SharedReg879_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_31_cast <= SharedReg879_out;
SharedReg110_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_32_cast <= SharedReg110_out;
SharedReg1107_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_33_cast <= SharedReg1107_out;
SharedReg114_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_34_cast <= SharedReg114_out;
SharedReg115_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_35_cast <= SharedReg115_out;
SharedReg1168_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_36_cast <= SharedReg1168_out;
SharedReg855_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_37_cast <= SharedReg855_out;
SharedReg642_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_38_cast <= SharedReg642_out;
SharedReg1160_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_39_cast <= SharedReg1160_out;
SharedReg290_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_40_cast <= SharedReg290_out;
SharedReg292_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_41_cast <= SharedReg292_out;
SharedReg1114_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_42_cast <= SharedReg1114_out;
SharedReg121_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_43_cast <= SharedReg121_out;
SharedReg861_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_44_cast <= SharedReg861_out;
SharedReg119_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_45_cast <= SharedReg119_out;
SharedReg646_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_46_cast <= SharedReg646_out;
SharedReg648_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_47_cast <= SharedReg648_out;
SharedReg1121_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_48_cast <= SharedReg1121_out;
SharedReg650_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_49_cast <= SharedReg650_out;
SharedReg1153_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_50_cast <= SharedReg1153_out;
SharedReg867_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_51_cast <= SharedReg867_out;
SharedReg296_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_52_cast <= SharedReg296_out;
SharedReg125_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_53_cast <= SharedReg125_out;
SharedReg651_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_54_cast <= SharedReg651_out;
SharedReg652_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_55_cast <= SharedReg652_out;
SharedReg124_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_56_cast <= SharedReg124_out;
SharedReg272_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_57_cast <= SharedReg272_out;
SharedReg125_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_58_cast <= SharedReg125_out;
SharedReg126_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_59_cast <= SharedReg126_out;
SharedReg269_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_60_cast <= SharedReg269_out;
SharedReg260_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_61_cast <= SharedReg260_out;
SharedReg640_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_62_cast <= SharedReg640_out;
SharedReg260_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_63_cast <= SharedReg260_out;
SharedReg234_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_64_cast <= SharedReg234_out;
   MUX_Product4_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg88_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg618_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg267_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg268_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg268_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg247_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg264_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg920_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg262_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1086_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg130_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg260_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg260_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg114_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg261_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg261_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg934_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg114_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1092_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg115_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg115_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg115_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg877_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg115_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg879_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg110_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1107_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg114_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg115_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1168_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg855_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg642_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1160_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg290_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg641_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg292_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1114_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg121_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg861_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg119_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg646_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg648_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1121_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg650_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1153_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg94_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg867_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg296_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg125_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg651_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg652_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg124_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg272_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg125_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg126_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg269_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg95_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg260_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg640_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg260_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg234_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg119_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg647_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg119_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product4_3_impl_1_out);

   Delay1No65_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_3_impl_1_out,
                 Y => Delay1No65_out);

Delay1No66_out_to_Product4_4_impl_parent_implementedSystem_port_0_cast <= Delay1No66_out;
Delay1No67_out_to_Product4_4_impl_parent_implementedSystem_port_1_cast <= Delay1No67_out;
   Product4_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_4_impl_out,
                 X => Delay1No66_out_to_Product4_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No67_out_to_Product4_4_impl_parent_implementedSystem_port_1_cast);

SharedReg1048_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1048_out;
SharedReg1049_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1049_out;
SharedReg1099_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1099_out;
SharedReg1051_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1051_out;
SharedReg1052_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1052_out;
SharedReg1019_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1019_out;
SharedReg1020_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1020_out;
SharedReg1021_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1021_out;
SharedReg1022_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1022_out;
SharedReg1023_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1023_out;
SharedReg1111_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1111_out;
SharedReg1024_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1024_out;
SharedReg1025_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1025_out;
SharedReg1113_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1113_out;
SharedReg1076_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1076_out;
SharedReg1027_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1027_out;
SharedReg1028_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1028_out;
SharedReg1029_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1029_out;
SharedReg1030_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1030_out;
SharedReg1031_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1031_out;
SharedReg1080_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1080_out;
SharedReg1032_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1032_out;
SharedReg1033_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1033_out;
SharedReg1034_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1034_out;
SharedReg1035_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1035_out;
SharedReg1085_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1085_out;
SharedReg125_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg125_out;
SharedReg1054_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1054_out;
SharedReg1038_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1038_out;
SharedReg1039_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1039_out;
SharedReg1040_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1040_out;
SharedReg1041_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1041_out;
SharedReg1130_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1130_out;
SharedReg1042_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1042_out;
SharedReg139_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_35_cast <= SharedReg139_out;
SharedReg1043_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1043_out;
SharedReg1044_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1044_out;
SharedReg1045_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1045_out;
SharedReg1104_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1104_out;
SharedReg1055_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1055_out;
SharedReg1056_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1056_out;
SharedReg679_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_42_cast <= SharedReg679_out;
SharedReg1057_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1057_out;
SharedReg1003_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1003_out;
SharedReg661_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_45_cast <= SharedReg661_out;
SharedReg1108_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1108_out;
SharedReg1154_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1154_out;
SharedReg858_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_48_cast <= SharedReg858_out;
SharedReg1007_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1007_out;
SharedReg1008_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1008_out;
SharedReg860_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_51_cast <= SharedReg860_out;
SharedReg1010_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1010_out;
SharedReg1150_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1150_out;
SharedReg1011_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1011_out;
SharedReg1123_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1123_out;
SharedReg1124_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1124_out;
SharedReg862_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_57_cast <= SharedReg862_out;
SharedReg1120_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1120_out;
SharedReg696_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_59_cast <= SharedReg696_out;
SharedReg1151_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1151_out;
SharedReg1016_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1016_out;
SharedReg1068_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1068_out;
SharedReg1161_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1161_out;
SharedReg1155_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1155_out;
   MUX_Product4_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1048_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1049_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1111_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1024_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1025_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1113_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1076_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1027_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1028_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1029_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1030_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1031_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1099_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1080_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1032_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1033_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1034_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1035_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1085_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg125_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1054_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1038_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1039_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1051_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1040_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1041_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1130_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1042_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg139_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1043_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1044_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1045_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1104_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1055_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1052_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1056_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg679_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1057_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1003_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg661_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1108_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1154_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg858_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1007_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1008_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1019_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg860_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1010_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1150_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1011_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1123_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1124_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg862_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1120_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg696_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1151_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1020_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1016_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1068_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1161_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1155_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1021_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1022_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1023_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product4_4_impl_0_out);

   Delay1No66_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_4_impl_0_out,
                 Y => Delay1No66_out);

SharedReg149_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg149_out;
SharedReg297_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg297_out;
SharedReg150_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg150_out;
SharedReg151_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg151_out;
SharedReg122_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg122_out;
SharedReg285_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg285_out;
SharedReg661_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg661_out;
SharedReg285_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg285_out;
SharedReg260_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg260_out;
SharedReg114_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg114_out;
SharedReg641_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg641_out;
SharedReg285_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg285_out;
SharedReg140_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg140_out;
SharedReg662_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg662_out;
SharedReg120_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg120_out;
SharedReg121_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg121_out;
SharedReg143_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg143_out;
SharedReg668_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg668_out;
SharedReg143_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg143_out;
SharedReg292_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg292_out;
SharedReg293_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg293_out;
SharedReg293_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg293_out;
SharedReg273_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg273_out;
SharedReg289_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg289_out;
SharedReg945_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg945_out;
SharedReg287_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg287_out;
SharedReg1086_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1086_out;
SharedReg305_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg305_out;
SharedReg285_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_29_cast <= SharedReg285_out;
SharedReg139_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_30_cast <= SharedReg139_out;
SharedReg286_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_31_cast <= SharedReg286_out;
SharedReg286_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_32_cast <= SharedReg286_out;
SharedReg858_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_33_cast <= SharedReg858_out;
SharedReg139_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_34_cast <= SharedReg139_out;
SharedReg1092_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_35_cast <= SharedReg1092_out;
SharedReg140_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_36_cast <= SharedReg140_out;
SharedReg140_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_37_cast <= SharedReg140_out;
SharedReg140_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_38_cast <= SharedReg140_out;
SharedReg680_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_39_cast <= SharedReg680_out;
SharedReg682_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_40_cast <= SharedReg682_out;
SharedReg280_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_41_cast <= SharedReg280_out;
SharedReg1107_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_42_cast <= SharedReg1107_out;
SharedReg139_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_43_cast <= SharedReg139_out;
SharedReg140_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_44_cast <= SharedReg140_out;
SharedReg1168_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_45_cast <= SharedReg1168_out;
SharedReg855_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_46_cast <= SharedReg855_out;
SharedReg857_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_47_cast <= SharedReg857_out;
SharedReg1160_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_48_cast <= SharedReg1160_out;
SharedReg315_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_49_cast <= SharedReg315_out;
SharedReg316_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_50_cast <= SharedReg316_out;
SharedReg1114_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_51_cast <= SharedReg1114_out;
SharedReg145_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_52_cast <= SharedReg145_out;
SharedReg667_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_53_cast <= SharedReg667_out;
SharedReg143_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_54_cast <= SharedReg143_out;
SharedReg667_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_55_cast <= SharedReg667_out;
SharedReg669_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_56_cast <= SharedReg669_out;
SharedReg1121_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1121_out;
SharedReg866_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_58_cast <= SharedReg866_out;
SharedReg1153_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_59_cast <= SharedReg1153_out;
SharedReg697_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_60_cast <= SharedReg697_out;
SharedReg319_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_61_cast <= SharedReg319_out;
SharedReg150_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_62_cast <= SharedReg150_out;
SharedReg674_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_63_cast <= SharedReg674_out;
SharedReg675_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_64_cast <= SharedReg675_out;
   MUX_Product4_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg149_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg297_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg641_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg285_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg140_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg662_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg120_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg121_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg143_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg668_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg143_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg292_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg150_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg293_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg293_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg273_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg289_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg945_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg287_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1086_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg305_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg285_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg139_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg151_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg286_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg286_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg858_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg139_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1092_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg140_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg140_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg140_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg680_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg682_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg122_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg280_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1107_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg139_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg140_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1168_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg855_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg857_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1160_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg315_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg316_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg285_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1114_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg145_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg667_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg143_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg667_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg669_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1121_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg866_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1153_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg697_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg661_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg319_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg150_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg674_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg675_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg285_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg260_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg114_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product4_4_impl_1_out);

   Delay1No67_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_4_impl_1_out,
                 Y => Delay1No67_out);

Delay1No68_out_to_Product4_5_impl_parent_implementedSystem_port_0_cast <= Delay1No68_out;
Delay1No69_out_to_Product4_5_impl_parent_implementedSystem_port_1_cast <= Delay1No69_out;
   Product4_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_5_impl_out,
                 X => Delay1No68_out_to_Product4_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No69_out_to_Product4_5_impl_parent_implementedSystem_port_1_cast);

SharedReg1124_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1124_out;
SharedReg692_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg692_out;
SharedReg1120_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1120_out;
SharedReg892_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg892_out;
SharedReg1151_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1151_out;
SharedReg1016_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1016_out;
SharedReg1068_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1068_out;
SharedReg1161_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1161_out;
SharedReg1155_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1155_out;
SharedReg1048_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1048_out;
SharedReg1049_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1049_out;
SharedReg1099_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1099_out;
SharedReg1051_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1051_out;
SharedReg1052_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1052_out;
SharedReg1019_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1019_out;
SharedReg1020_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1020_out;
SharedReg1021_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1021_out;
SharedReg1022_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1022_out;
SharedReg1023_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1023_out;
SharedReg1111_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1111_out;
SharedReg1024_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1024_out;
SharedReg1025_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1025_out;
SharedReg1113_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1113_out;
SharedReg1076_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1076_out;
SharedReg1027_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1027_out;
SharedReg1028_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1028_out;
SharedReg1029_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1029_out;
SharedReg1030_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1030_out;
SharedReg1031_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1031_out;
SharedReg1080_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1080_out;
SharedReg1032_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1032_out;
SharedReg1033_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1033_out;
SharedReg1034_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1034_out;
SharedReg1035_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1035_out;
SharedReg1085_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1085_out;
SharedReg150_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_36_cast <= SharedReg150_out;
SharedReg1054_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1054_out;
SharedReg1038_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1038_out;
SharedReg1039_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1039_out;
SharedReg1040_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1040_out;
SharedReg1041_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1041_out;
SharedReg1130_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1130_out;
SharedReg1042_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1042_out;
SharedReg163_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_44_cast <= SharedReg163_out;
SharedReg1043_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1043_out;
SharedReg1044_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1044_out;
SharedReg1045_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1045_out;
SharedReg1104_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1104_out;
SharedReg1055_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1055_out;
SharedReg1056_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1056_out;
SharedReg723_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_51_cast <= SharedReg723_out;
SharedReg1057_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1057_out;
SharedReg1003_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1003_out;
SharedReg707_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_54_cast <= SharedReg707_out;
SharedReg1108_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1108_out;
SharedReg1154_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1154_out;
SharedReg688_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_57_cast <= SharedReg688_out;
SharedReg1007_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1007_out;
SharedReg1008_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1008_out;
SharedReg690_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_60_cast <= SharedReg690_out;
SharedReg1010_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1010_out;
SharedReg1150_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1150_out;
SharedReg1011_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1011_out;
SharedReg1123_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1123_out;
   MUX_Product4_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1124_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg692_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1049_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1099_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1051_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1052_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1019_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1020_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1021_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1022_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1023_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1111_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1120_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1024_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1025_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1113_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1076_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1027_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1028_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1029_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1030_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1031_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1080_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg892_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1032_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1033_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1034_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1035_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1085_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg150_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1054_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1038_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1039_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1040_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1151_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1041_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1130_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1042_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg163_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1043_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1044_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1045_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1104_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1055_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1056_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1016_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg723_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1057_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1003_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg707_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1108_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1154_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg688_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1007_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1008_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg690_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1068_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1010_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1150_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1011_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1123_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1161_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1155_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1048_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product4_5_impl_0_out);

   Delay1No68_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_5_impl_0_out,
                 Y => Delay1No68_out);

SharedReg715_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg715_out;
SharedReg1121_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1121_out;
SharedReg672_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg672_out;
SharedReg1153_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1153_out;
SharedReg893_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg893_out;
SharedReg197_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg197_out;
SharedReg175_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg175_out;
SharedReg718_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg718_out;
SharedReg719_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg719_out;
SharedReg320_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg320_out;
SharedReg149_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg149_out;
SharedReg321_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg321_out;
SharedReg322_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg322_out;
SharedReg294_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_14_cast <= SharedReg294_out;
SharedReg310_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_15_cast <= SharedReg310_out;
SharedReg707_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_16_cast <= SharedReg707_out;
SharedReg310_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_17_cast <= SharedReg310_out;
SharedReg285_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_18_cast <= SharedReg285_out;
SharedReg139_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_19_cast <= SharedReg139_out;
SharedReg662_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_20_cast <= SharedReg662_out;
SharedReg310_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_21_cast <= SharedReg310_out;
SharedReg164_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_22_cast <= SharedReg164_out;
SharedReg708_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_23_cast <= SharedReg708_out;
SharedReg144_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_24_cast <= SharedReg144_out;
SharedReg145_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_25_cast <= SharedReg145_out;
SharedReg169_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_26_cast <= SharedReg169_out;
SharedReg714_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_27_cast <= SharedReg714_out;
SharedReg169_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_28_cast <= SharedReg169_out;
SharedReg316_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_29_cast <= SharedReg316_out;
SharedReg317_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_30_cast <= SharedReg317_out;
SharedReg317_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_31_cast <= SharedReg317_out;
SharedReg298_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_32_cast <= SharedReg298_out;
SharedReg314_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_33_cast <= SharedReg314_out;
SharedReg870_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_34_cast <= SharedReg870_out;
SharedReg141_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_35_cast <= SharedReg141_out;
SharedReg1086_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_36_cast <= SharedReg1086_out;
SharedReg327_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_37_cast <= SharedReg327_out;
SharedReg310_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_38_cast <= SharedReg310_out;
SharedReg163_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_39_cast <= SharedReg163_out;
SharedReg311_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_40_cast <= SharedReg311_out;
SharedReg311_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_41_cast <= SharedReg311_out;
SharedReg688_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_42_cast <= SharedReg688_out;
SharedReg163_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_43_cast <= SharedReg163_out;
SharedReg1092_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_44_cast <= SharedReg1092_out;
SharedReg164_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_45_cast <= SharedReg164_out;
SharedReg311_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_46_cast <= SharedReg311_out;
SharedReg140_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_47_cast <= SharedReg140_out;
SharedReg724_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_48_cast <= SharedReg724_out;
SharedReg726_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_49_cast <= SharedReg726_out;
SharedReg306_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_50_cast <= SharedReg306_out;
SharedReg1107_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_51_cast <= SharedReg1107_out;
SharedReg163_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_52_cast <= SharedReg163_out;
SharedReg164_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_53_cast <= SharedReg164_out;
SharedReg1168_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_54_cast <= SharedReg1168_out;
SharedReg685_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_55_cast <= SharedReg685_out;
SharedReg687_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_56_cast <= SharedReg687_out;
SharedReg1160_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1160_out;
SharedReg191_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_58_cast <= SharedReg191_out;
SharedReg193_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_59_cast <= SharedReg193_out;
SharedReg1114_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_60_cast <= SharedReg1114_out;
SharedReg171_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_61_cast <= SharedReg171_out;
SharedReg691_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_62_cast <= SharedReg691_out;
SharedReg169_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_63_cast <= SharedReg169_out;
SharedReg713_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_64_cast <= SharedReg713_out;
   MUX_Product4_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg715_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1121_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg149_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg321_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg322_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg294_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg310_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg707_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg310_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg285_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg139_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg662_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg672_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg310_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg164_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg708_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg144_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg145_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg169_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg714_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg169_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg316_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg317_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1153_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg317_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg298_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg314_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg870_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg141_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1086_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg327_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg310_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg163_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg311_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg893_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg311_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg688_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg163_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1092_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg164_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg311_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg140_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg724_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg726_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg306_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg197_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1107_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg163_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg164_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1168_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg685_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg687_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1160_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg191_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg193_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1114_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg175_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg171_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg691_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg169_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg713_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg718_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg719_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg320_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product4_5_impl_1_out);

   Delay1No69_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_5_impl_1_out,
                 Y => Delay1No69_out);

Delay1No70_out_to_Product4_6_impl_parent_implementedSystem_port_0_cast <= Delay1No70_out;
Delay1No71_out_to_Product4_6_impl_parent_implementedSystem_port_1_cast <= Delay1No71_out;
   Product4_6_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_6_impl_out,
                 X => Delay1No70_out_to_Product4_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No71_out_to_Product4_6_impl_parent_implementedSystem_port_1_cast);

SharedReg1108_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1108_out;
SharedReg1154_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1154_out;
SharedReg688_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg688_out;
SharedReg1007_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1007_out;
SharedReg1008_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1008_out;
SharedReg712_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg712_out;
SharedReg1010_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1010_out;
SharedReg1150_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1150_out;
SharedReg1011_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1011_out;
SharedReg1123_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1123_out;
SharedReg1124_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1124_out;
SharedReg714_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg714_out;
SharedReg1120_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1120_out;
SharedReg994_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_14_cast <= SharedReg994_out;
SharedReg1151_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1151_out;
SharedReg1016_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1016_out;
SharedReg1068_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1068_out;
SharedReg1161_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1161_out;
SharedReg1155_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1155_out;
SharedReg1048_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1048_out;
SharedReg1049_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1049_out;
SharedReg1099_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1099_out;
SharedReg1051_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1051_out;
SharedReg1052_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1052_out;
SharedReg1019_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1019_out;
SharedReg1020_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1020_out;
SharedReg1021_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1021_out;
SharedReg1022_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1022_out;
SharedReg1023_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1023_out;
SharedReg1111_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1111_out;
SharedReg1024_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1024_out;
SharedReg1025_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1025_out;
SharedReg1113_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1113_out;
SharedReg1076_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1076_out;
SharedReg1027_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1027_out;
SharedReg1028_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1028_out;
SharedReg1029_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1029_out;
SharedReg1030_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1030_out;
SharedReg1031_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1031_out;
SharedReg1080_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1080_out;
SharedReg1032_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1032_out;
SharedReg1033_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1033_out;
SharedReg1034_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1034_out;
SharedReg1035_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1035_out;
SharedReg1085_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1085_out;
SharedReg175_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_46_cast <= SharedReg175_out;
SharedReg1054_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1054_out;
SharedReg1038_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1038_out;
SharedReg1039_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1039_out;
SharedReg1040_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1040_out;
SharedReg1041_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1041_out;
SharedReg1130_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1130_out;
SharedReg1042_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1042_out;
SharedReg186_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_54_cast <= SharedReg186_out;
SharedReg1043_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1043_out;
SharedReg1044_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1044_out;
SharedReg1045_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1045_out;
SharedReg1104_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1104_out;
SharedReg1055_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1055_out;
SharedReg1056_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1056_out;
SharedReg999_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_61_cast <= SharedReg999_out;
SharedReg1057_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1057_out;
SharedReg1003_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1003_out;
SharedReg707_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_64_cast <= SharedReg707_out;
   MUX_Product4_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1108_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1154_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1124_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg714_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1120_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg994_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1151_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1016_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1068_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1161_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1155_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1048_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg688_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1049_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1099_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1051_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1052_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1019_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1020_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1021_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1022_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1023_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1111_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1007_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1024_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1025_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1113_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1076_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1027_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1028_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1029_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1030_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1031_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1080_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1008_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1032_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1033_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1034_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1035_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1085_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg175_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1054_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1038_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1039_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1040_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg712_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1041_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1130_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1042_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg186_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1043_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1044_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1045_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1104_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1055_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1056_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1010_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg999_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1057_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1003_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg707_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1150_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1011_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1123_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product4_6_impl_0_out);

   Delay1No70_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_6_impl_0_out,
                 Y => Delay1No70_out);

SharedReg707_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg707_out;
SharedReg687_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg687_out;
SharedReg1160_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1160_out;
SharedReg191_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg191_out;
SharedReg339_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg339_out;
SharedReg1114_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1114_out;
SharedReg171_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg171_out;
SharedReg989_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg989_out;
SharedReg192_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg192_out;
SharedReg713_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg713_out;
SharedReg890_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg890_out;
SharedReg1121_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1121_out;
SharedReg892_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_13_cast <= SharedReg892_out;
SharedReg1153_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1153_out;
SharedReg995_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_15_cast <= SharedReg995_out;
SharedReg173_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_16_cast <= SharedReg173_out;
SharedReg199_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_17_cast <= SharedReg199_out;
SharedReg894_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_18_cast <= SharedReg894_out;
SharedReg895_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_19_cast <= SharedReg895_out;
SharedReg174_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_20_cast <= SharedReg174_out;
SharedReg320_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_21_cast <= SharedReg320_out;
SharedReg175_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_22_cast <= SharedReg175_out;
SharedReg176_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_23_cast <= SharedReg176_out;
SharedReg195_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_24_cast <= SharedReg195_out;
SharedReg186_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_25_cast <= SharedReg186_out;
SharedReg882_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_26_cast <= SharedReg882_out;
SharedReg163_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_27_cast <= SharedReg163_out;
SharedReg310_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_28_cast <= SharedReg310_out;
SharedReg332_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_29_cast <= SharedReg332_out;
SharedReg984_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_30_cast <= SharedReg984_out;
SharedReg186_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_31_cast <= SharedReg186_out;
SharedReg333_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_32_cast <= SharedReg333_out;
SharedReg708_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_33_cast <= SharedReg708_out;
SharedReg316_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_34_cast <= SharedReg316_out;
SharedReg317_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_35_cast <= SharedReg317_out;
SharedReg338_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_36_cast <= SharedReg338_out;
SharedReg990_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_37_cast <= SharedReg990_out;
SharedReg192_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_38_cast <= SharedReg192_out;
SharedReg170_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_39_cast <= SharedReg170_out;
SharedReg171_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_40_cast <= SharedReg171_out;
SharedReg194_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_41_cast <= SharedReg194_out;
SharedReg199_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_42_cast <= SharedReg199_out;
SharedReg190_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_43_cast <= SharedReg190_out;
SharedReg896_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_44_cast <= SharedReg896_out;
SharedReg188_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_45_cast <= SharedReg188_out;
SharedReg1086_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_46_cast <= SharedReg1086_out;
SharedReg178_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_47_cast <= SharedReg178_out;
SharedReg186_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_48_cast <= SharedReg186_out;
SharedReg332_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_49_cast <= SharedReg332_out;
SharedReg187_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_50_cast <= SharedReg187_out;
SharedReg187_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_51_cast <= SharedReg187_out;
SharedReg885_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_52_cast <= SharedReg885_out;
SharedReg332_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_53_cast <= SharedReg332_out;
SharedReg1092_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_54_cast <= SharedReg1092_out;
SharedReg187_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_55_cast <= SharedReg187_out;
SharedReg164_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_56_cast <= SharedReg164_out;
SharedReg164_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_57_cast <= SharedReg164_out;
SharedReg901_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_58_cast <= SharedReg901_out;
SharedReg1000_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_59_cast <= SharedReg1000_out;
SharedReg205_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_60_cast <= SharedReg205_out;
SharedReg1107_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_61_cast <= SharedReg1107_out;
SharedReg186_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_62_cast <= SharedReg186_out;
SharedReg187_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_63_cast <= SharedReg187_out;
SharedReg1168_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_64_cast <= SharedReg1168_out;
   MUX_Product4_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg707_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg687_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg890_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1121_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg892_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1153_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg995_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg173_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg199_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg894_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg895_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg174_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1160_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg320_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg175_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg176_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg195_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg186_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg882_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg163_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg310_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg332_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg984_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg191_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg186_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg333_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg708_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg316_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg317_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg338_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg990_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg192_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg170_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg171_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg339_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg194_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg199_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg190_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg896_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg188_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1086_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg178_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg186_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg332_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg187_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1114_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg187_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg885_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg332_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1092_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg187_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg164_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg164_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg901_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1000_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg205_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg171_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1107_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg186_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg187_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1168_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg989_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg192_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg713_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product4_6_impl_1_out);

   Delay1No71_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_6_impl_1_out,
                 Y => Delay1No71_out);

Delay1No72_out_to_Product31_0_impl_parent_implementedSystem_port_0_cast <= Delay1No72_out;
Delay1No73_out_to_Product31_0_impl_parent_implementedSystem_port_1_cast <= Delay1No73_out;
   Product31_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product31_0_impl_out,
                 X => Delay1No72_out_to_Product31_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No73_out_to_Product31_0_impl_parent_implementedSystem_port_1_cast);

SharedReg37_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg37_out;
SharedReg1094_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1094_out;
SharedReg1135_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1135_out;
SharedReg1105_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1105_out;
SharedReg57_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg57_out;
SharedReg1046_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1046_out;
SharedReg1057_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1057_out;
SharedReg1170_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1170_out;
SharedReg1004_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1004_out;
SharedReg1166_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1166_out;
SharedReg1006_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1006_out;
SharedReg1171_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1171_out;
SharedReg1060_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1060_out;
SharedReg215_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg215_out;
SharedReg213_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg213_out;
SharedReg1115_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1115_out;
SharedReg1152_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1152_out;
SharedReg1063_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1063_out;
SharedReg1136_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1136_out;
SharedReg575_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg575_out;
SharedReg1013_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1013_out;
SharedReg1120_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1120_out;
SharedReg1014_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1014_out;
SharedReg1015_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1015_out;
SharedReg219_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg219_out;
SharedReg1017_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1017_out;
SharedReg1018_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1018_out;
SharedReg1047_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1047_out;
SharedReg48_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_29_cast <= SharedReg48_out;
SharedReg1049_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1049_out;
SharedReg1050_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1050_out;
SharedReg1051_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1051_out;
SharedReg45_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_33_cast <= SharedReg45_out;
SharedReg36_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_34_cast <= SharedReg36_out;
SharedReg957_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_35_cast <= SharedReg957_out;
SharedReg1156_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1156_out;
SharedReg1072_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1072_out;
SharedReg208_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_38_cast <= SharedReg208_out;
SharedReg958_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_39_cast <= SharedReg958_out;
SharedReg1074_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1074_out;
SharedReg209_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_41_cast <= SharedReg209_out;
SharedReg958_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_42_cast <= SharedReg958_out;
SharedReg215_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_43_cast <= SharedReg215_out;
SharedReg1158_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1158_out;
SharedReg1077_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1077_out;
SharedReg1029_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1029_out;
SharedReg214_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_47_cast <= SharedReg214_out;
SharedReg1159_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1159_out;
SharedReg1125_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1125_out;
SharedReg1081_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1081_out;
SharedReg1082_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1082_out;
SharedReg40_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_52_cast <= SharedReg40_out;
SharedReg1084_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1084_out;
SharedReg1036_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1036_out;
SharedReg1037_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1037_out;
SharedReg1103_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1103_out;
SharedReg36_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_57_cast <= SharedReg36_out;
SharedReg208_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_58_cast <= SharedReg208_out;
SharedReg1089_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1089_out;
SharedReg1090_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1090_out;
SharedReg1145_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1145_out;
SharedReg1091_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1091_out;
SharedReg1132_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1132_out;
SharedReg1133_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1133_out;
   MUX_Product31_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg37_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1094_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1006_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1171_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1060_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg215_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg213_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1115_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1152_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1063_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1136_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg575_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1135_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1013_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1120_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1014_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1015_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg219_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1017_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1018_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1047_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg48_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1049_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1105_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1050_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1051_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg45_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg36_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg957_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1156_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1072_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg208_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg958_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1074_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg57_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg209_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg958_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg215_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1158_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1077_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1029_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg214_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1159_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1125_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1081_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1046_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1082_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg40_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1084_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1036_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1037_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1103_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg36_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg208_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1089_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1090_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1057_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1145_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1091_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1132_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1133_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1170_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1004_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1166_out_to_MUX_Product31_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product31_0_impl_0_out);

   Delay1No72_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_0_impl_0_out,
                 Y => Delay1No72_out);

SharedReg1093_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1093_out;
SharedReg37_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg37_out;
SharedReg569_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg569_out;
SharedReg980_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg980_out;
SharedReg1106_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1106_out;
SharedReg36_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg36_out;
SharedReg567_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg567_out;
SharedReg567_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg567_out;
SharedReg36_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg36_out;
SharedReg958_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg958_out;
SharedReg37_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg37_out;
SharedReg571_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg571_out;
SharedReg41_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg41_out;
SharedReg1061_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1061_out;
SharedReg1062_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1062_out;
SharedReg573_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg573_out;
SharedReg963_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg963_out;
SharedReg213_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg213_out;
SharedReg573_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg573_out;
SharedReg1137_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1137_out;
SharedReg46_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg46_out;
SharedReg575_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg575_out;
SharedReg218_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg218_out;
SharedReg220_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg220_out;
SharedReg1067_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1067_out;
SharedReg223_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg223_out;
SharedReg49_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg49_out;
SharedReg577_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg577_out;
SharedReg1097_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_29_cast <= SharedReg1097_out;
SharedReg578_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_30_cast <= SharedReg578_out;
SharedReg971_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_31_cast <= SharedReg971_out;
SharedReg971_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_32_cast <= SharedReg971_out;
SharedReg1101_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_33_cast <= SharedReg1101_out;
SharedReg1070_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_34_cast <= SharedReg1070_out;
SharedReg1071_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_35_cast <= SharedReg1071_out;
SharedReg567_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_36_cast <= SharedReg567_out;
SharedReg36_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_37_cast <= SharedReg36_out;
SharedReg1073_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_38_cast <= SharedReg1073_out;
SharedReg1117_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_39_cast <= SharedReg1117_out;
SharedReg36_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_40_cast <= SharedReg36_out;
SharedReg1075_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_41_cast <= SharedReg1075_out;
SharedReg1119_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_42_cast <= SharedReg1119_out;
SharedReg1076_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_43_cast <= SharedReg1076_out;
SharedReg965_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_44_cast <= SharedReg965_out;
SharedReg214_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_45_cast <= SharedReg214_out;
SharedReg573_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_46_cast <= SharedReg573_out;
SharedReg1079_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_47_cast <= SharedReg1079_out;
SharedReg574_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_48_cast <= SharedReg574_out;
SharedReg574_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_49_cast <= SharedReg574_out;
SharedReg216_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_50_cast <= SharedReg216_out;
SharedReg49_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_51_cast <= SharedReg49_out;
SharedReg1083_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_52_cast <= SharedReg1083_out;
SharedReg580_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_53_cast <= SharedReg580_out;
SharedReg38_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_54_cast <= SharedReg38_out;
SharedReg49_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_55_cast <= SharedReg49_out;
SharedReg56_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_56_cast <= SharedReg56_out;
SharedReg1087_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1087_out;
SharedReg1088_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_58_cast <= SharedReg1088_out;
SharedReg37_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_59_cast <= SharedReg37_out;
SharedReg37_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_60_cast <= SharedReg37_out;
SharedReg570_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_61_cast <= SharedReg570_out;
SharedReg36_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_62_cast <= SharedReg36_out;
SharedReg568_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_63_cast <= SharedReg568_out;
SharedReg568_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_64_cast <= SharedReg568_out;
   MUX_Product31_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1093_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg37_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg37_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg571_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg41_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1061_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1062_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg573_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg963_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg213_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg573_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1137_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg569_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg46_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg575_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg218_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg220_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1067_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg223_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg49_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg577_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1097_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg578_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg980_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg971_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg971_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1101_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1070_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1071_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg567_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg36_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1073_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1117_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg36_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1106_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1075_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1119_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1076_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg965_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg214_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg573_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1079_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg574_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg574_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg216_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg36_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg49_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1083_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg580_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg38_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg49_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg56_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1087_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1088_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg37_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg37_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg567_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg570_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg36_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg568_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg568_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg567_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg36_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg958_out_to_MUX_Product31_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product31_0_impl_1_out);

   Delay1No73_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_0_impl_1_out,
                 Y => Delay1No73_out);

Delay1No74_out_to_Product31_1_impl_parent_implementedSystem_port_0_cast <= Delay1No74_out;
Delay1No75_out_to_Product31_1_impl_parent_implementedSystem_port_1_cast <= Delay1No75_out;
   Product31_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product31_1_impl_out,
                 X => Delay1No74_out_to_Product31_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No75_out_to_Product31_1_impl_parent_implementedSystem_port_1_cast);

SharedReg1103_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1103_out;
SharedReg208_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg208_out;
SharedReg62_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg62_out;
SharedReg1089_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1089_out;
SharedReg1090_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1090_out;
SharedReg1145_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1145_out;
SharedReg1091_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1091_out;
SharedReg1132_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1132_out;
SharedReg1133_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1133_out;
SharedReg63_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg63_out;
SharedReg1094_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1094_out;
SharedReg1135_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1135_out;
SharedReg1105_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1105_out;
SharedReg83_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg83_out;
SharedReg1046_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1046_out;
SharedReg1057_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1057_out;
SharedReg1170_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1170_out;
SharedReg1004_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1004_out;
SharedReg1166_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1166_out;
SharedReg1006_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1006_out;
SharedReg1171_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1171_out;
SharedReg1060_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1060_out;
SharedReg241_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg241_out;
SharedReg239_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg239_out;
SharedReg1115_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1115_out;
SharedReg1152_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1152_out;
SharedReg1063_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1063_out;
SharedReg1136_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1136_out;
SharedReg601_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_29_cast <= SharedReg601_out;
SharedReg1013_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1013_out;
SharedReg1120_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1120_out;
SharedReg1014_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1014_out;
SharedReg1015_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1015_out;
SharedReg245_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_34_cast <= SharedReg245_out;
SharedReg1017_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1017_out;
SharedReg1018_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1018_out;
SharedReg1047_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1047_out;
SharedReg74_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_38_cast <= SharedReg74_out;
SharedReg1049_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1049_out;
SharedReg1050_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1050_out;
SharedReg1051_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1051_out;
SharedReg217_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_42_cast <= SharedReg217_out;
SharedReg62_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_43_cast <= SharedReg62_out;
SharedReg906_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_44_cast <= SharedReg906_out;
SharedReg1156_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1156_out;
SharedReg1072_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1072_out;
SharedReg62_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_47_cast <= SharedReg62_out;
SharedReg594_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_48_cast <= SharedReg594_out;
SharedReg1074_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1074_out;
SharedReg235_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_50_cast <= SharedReg235_out;
SharedReg907_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_51_cast <= SharedReg907_out;
SharedReg69_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_52_cast <= SharedReg69_out;
SharedReg1158_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1158_out;
SharedReg1077_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1077_out;
SharedReg1029_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1029_out;
SharedReg240_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_56_cast <= SharedReg240_out;
SharedReg1159_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1159_out;
SharedReg1125_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1125_out;
SharedReg1081_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1081_out;
SharedReg1082_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1082_out;
SharedReg66_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_61_cast <= SharedReg66_out;
SharedReg1084_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1084_out;
SharedReg1036_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1036_out;
SharedReg1037_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1037_out;
   MUX_Product31_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1103_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg208_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1094_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1135_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1105_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg83_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1046_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1057_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1170_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1004_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1166_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1006_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg62_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1171_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1060_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg241_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg239_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1115_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1152_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1063_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1136_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg601_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1013_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1089_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1120_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1014_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1015_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg245_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1017_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1018_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1047_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg74_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1049_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1050_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1090_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1051_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg217_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg62_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg906_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1156_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1072_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg62_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg594_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1074_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg235_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1145_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg907_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg69_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1158_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1077_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1029_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg240_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1159_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1125_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1081_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1082_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1091_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg66_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1084_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1036_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1037_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1132_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1133_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg63_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product31_1_impl_0_out);

   Delay1No74_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_1_impl_0_out,
                 Y => Delay1No74_out);

SharedReg80_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg80_out;
SharedReg1087_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1087_out;
SharedReg1088_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1088_out;
SharedReg209_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg209_out;
SharedReg209_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg209_out;
SharedReg960_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg960_out;
SharedReg62_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg62_out;
SharedReg594_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg594_out;
SharedReg594_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg594_out;
SharedReg1093_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1093_out;
SharedReg63_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg63_out;
SharedReg595_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg595_out;
SharedReg928_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg928_out;
SharedReg1106_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1106_out;
SharedReg62_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg62_out;
SharedReg593_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg593_out;
SharedReg593_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg593_out;
SharedReg62_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg62_out;
SharedReg907_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg907_out;
SharedReg63_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg63_out;
SharedReg597_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg597_out;
SharedReg67_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg67_out;
SharedReg1061_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1061_out;
SharedReg1062_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1062_out;
SharedReg599_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg599_out;
SharedReg912_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg912_out;
SharedReg239_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg239_out;
SharedReg599_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg599_out;
SharedReg1137_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_29_cast <= SharedReg1137_out;
SharedReg72_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_30_cast <= SharedReg72_out;
SharedReg965_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_31_cast <= SharedReg965_out;
SharedReg244_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_32_cast <= SharedReg244_out;
SharedReg246_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_33_cast <= SharedReg246_out;
SharedReg1067_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_34_cast <= SharedReg1067_out;
SharedReg249_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_35_cast <= SharedReg249_out;
SharedReg75_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_36_cast <= SharedReg75_out;
SharedReg603_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_37_cast <= SharedReg603_out;
SharedReg1097_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_38_cast <= SharedReg1097_out;
SharedReg604_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_39_cast <= SharedReg604_out;
SharedReg919_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_40_cast <= SharedReg919_out;
SharedReg919_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_41_cast <= SharedReg919_out;
SharedReg1101_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_42_cast <= SharedReg1101_out;
SharedReg1070_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_43_cast <= SharedReg1070_out;
SharedReg1071_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_44_cast <= SharedReg1071_out;
SharedReg957_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_45_cast <= SharedReg957_out;
SharedReg36_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_46_cast <= SharedReg36_out;
SharedReg1073_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_47_cast <= SharedReg1073_out;
SharedReg1117_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_48_cast <= SharedReg1117_out;
SharedReg62_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_49_cast <= SharedReg62_out;
SharedReg1075_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_50_cast <= SharedReg1075_out;
SharedReg1119_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_51_cast <= SharedReg1119_out;
SharedReg1076_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_52_cast <= SharedReg1076_out;
SharedReg601_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_53_cast <= SharedReg601_out;
SharedReg240_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_54_cast <= SharedReg240_out;
SharedReg599_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_55_cast <= SharedReg599_out;
SharedReg1079_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_56_cast <= SharedReg1079_out;
SharedReg600_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_57_cast <= SharedReg600_out;
SharedReg600_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_58_cast <= SharedReg600_out;
SharedReg242_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_59_cast <= SharedReg242_out;
SharedReg221_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_60_cast <= SharedReg221_out;
SharedReg1083_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_61_cast <= SharedReg1083_out;
SharedReg972_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_62_cast <= SharedReg972_out;
SharedReg210_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_63_cast <= SharedReg210_out;
SharedReg75_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_64_cast <= SharedReg75_out;
   MUX_Product31_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg80_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1087_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg63_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg595_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg928_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1106_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg62_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg593_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg593_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg62_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg907_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg63_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1088_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg597_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg67_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1061_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1062_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg599_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg912_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg239_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg599_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1137_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg72_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg209_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg965_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg244_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg246_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1067_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg249_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg75_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg603_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1097_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg604_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg919_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg209_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg919_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1101_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1070_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1071_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg957_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg36_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1073_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1117_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg62_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1075_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg960_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1119_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1076_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg601_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg240_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg599_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1079_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg600_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg600_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg242_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg221_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg62_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1083_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg972_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg210_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg75_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg594_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg594_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1093_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product31_1_impl_1_out);

   Delay1No75_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_1_impl_1_out,
                 Y => Delay1No75_out);

Delay1No76_out_to_Product31_2_impl_parent_implementedSystem_port_0_cast <= Delay1No76_out;
Delay1No77_out_to_Product31_2_impl_parent_implementedSystem_port_1_cast <= Delay1No77_out;
   Product31_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product31_2_impl_out,
                 X => Delay1No76_out_to_Product31_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No77_out_to_Product31_2_impl_parent_implementedSystem_port_1_cast);

SharedReg266_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg266_out;
SharedReg1159_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1159_out;
SharedReg1125_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1125_out;
SharedReg1081_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1081_out;
SharedReg1082_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1082_out;
SharedReg238_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg238_out;
SharedReg1084_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1084_out;
SharedReg1036_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1036_out;
SharedReg1037_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1037_out;
SharedReg1103_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1103_out;
SharedReg234_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg234_out;
SharedReg88_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg88_out;
SharedReg1089_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1089_out;
SharedReg1090_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1090_out;
SharedReg1145_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1145_out;
SharedReg1091_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1091_out;
SharedReg1132_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1132_out;
SharedReg1133_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1133_out;
SharedReg89_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg89_out;
SharedReg1094_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1094_out;
SharedReg1135_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1135_out;
SharedReg1105_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1105_out;
SharedReg255_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg255_out;
SharedReg1046_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1046_out;
SharedReg1057_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1057_out;
SharedReg1170_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1170_out;
SharedReg1004_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1004_out;
SharedReg1166_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1166_out;
SharedReg1006_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1006_out;
SharedReg1171_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1171_out;
SharedReg1060_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1060_out;
SharedReg267_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_32_cast <= SharedReg267_out;
SharedReg265_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_33_cast <= SharedReg265_out;
SharedReg1115_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1115_out;
SharedReg1152_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1152_out;
SharedReg1063_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1063_out;
SharedReg1136_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1136_out;
SharedReg625_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_38_cast <= SharedReg625_out;
SharedReg1013_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1013_out;
SharedReg1120_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1120_out;
SharedReg1014_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1014_out;
SharedReg1015_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1015_out;
SharedReg271_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_43_cast <= SharedReg271_out;
SharedReg1017_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1017_out;
SharedReg1018_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1018_out;
SharedReg1047_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1047_out;
SharedReg99_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_47_cast <= SharedReg99_out;
SharedReg1049_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1049_out;
SharedReg1050_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1050_out;
SharedReg1051_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1051_out;
SharedReg243_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_51_cast <= SharedReg243_out;
SharedReg88_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_52_cast <= SharedReg88_out;
SharedReg931_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_53_cast <= SharedReg931_out;
SharedReg1156_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1156_out;
SharedReg1072_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1072_out;
SharedReg234_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_56_cast <= SharedReg234_out;
SharedReg907_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_57_cast <= SharedReg907_out;
SharedReg1074_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1074_out;
SharedReg261_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_59_cast <= SharedReg261_out;
SharedReg932_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_60_cast <= SharedReg932_out;
SharedReg94_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_61_cast <= SharedReg94_out;
SharedReg1158_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1158_out;
SharedReg1077_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1077_out;
SharedReg1029_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1029_out;
   MUX_Product31_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg266_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1159_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg234_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg88_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1089_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1090_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1145_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1091_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1132_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1133_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg89_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1094_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1125_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1135_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1105_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg255_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1046_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1057_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1170_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1004_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1166_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1006_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1171_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1081_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1060_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg267_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg265_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1115_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1152_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1063_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1136_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg625_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1013_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1120_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1082_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1014_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1015_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg271_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1017_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1018_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1047_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg99_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1049_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1050_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1051_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg238_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg243_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg88_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg931_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1156_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1072_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg234_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg907_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1074_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg261_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg932_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1084_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg94_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1158_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1077_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1029_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1036_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1037_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1103_out_to_MUX_Product31_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product31_2_impl_0_out);

   Delay1No76_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_2_impl_0_out,
                 Y => Delay1No76_out);

SharedReg1079_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1079_out;
SharedReg624_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg624_out;
SharedReg913_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg913_out;
SharedReg95_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg95_out;
SharedReg75_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg75_out;
SharedReg1083_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1083_out;
SharedReg607_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg607_out;
SharedReg236_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg236_out;
SharedReg247_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg247_out;
SharedReg105_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg105_out;
SharedReg1087_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1087_out;
SharedReg1088_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1088_out;
SharedReg235_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg235_out;
SharedReg235_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg235_out;
SharedReg909_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg909_out;
SharedReg88_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg88_out;
SharedReg618_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg618_out;
SharedReg618_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg618_out;
SharedReg1093_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1093_out;
SharedReg89_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg89_out;
SharedReg619_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg619_out;
SharedReg954_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg954_out;
SharedReg1106_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1106_out;
SharedReg88_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg88_out;
SharedReg617_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg617_out;
SharedReg617_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg617_out;
SharedReg88_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg88_out;
SharedReg932_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg932_out;
SharedReg89_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_29_cast <= SharedReg89_out;
SharedReg621_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_30_cast <= SharedReg621_out;
SharedReg92_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_31_cast <= SharedReg92_out;
SharedReg1061_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_32_cast <= SharedReg1061_out;
SharedReg1062_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_33_cast <= SharedReg1062_out;
SharedReg623_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_34_cast <= SharedReg623_out;
SharedReg937_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_35_cast <= SharedReg937_out;
SharedReg265_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_36_cast <= SharedReg265_out;
SharedReg623_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_37_cast <= SharedReg623_out;
SharedReg1137_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_38_cast <= SharedReg1137_out;
SharedReg97_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_39_cast <= SharedReg97_out;
SharedReg914_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_40_cast <= SharedReg914_out;
SharedReg270_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_41_cast <= SharedReg270_out;
SharedReg272_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_42_cast <= SharedReg272_out;
SharedReg1067_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_43_cast <= SharedReg1067_out;
SharedReg275_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_44_cast <= SharedReg275_out;
SharedReg100_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_45_cast <= SharedReg100_out;
SharedReg628_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_46_cast <= SharedReg628_out;
SharedReg1097_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_47_cast <= SharedReg1097_out;
SharedReg629_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_48_cast <= SharedReg629_out;
SharedReg944_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_49_cast <= SharedReg944_out;
SharedReg944_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_50_cast <= SharedReg944_out;
SharedReg1101_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_51_cast <= SharedReg1101_out;
SharedReg1070_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_52_cast <= SharedReg1070_out;
SharedReg1071_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_53_cast <= SharedReg1071_out;
SharedReg906_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_54_cast <= SharedReg906_out;
SharedReg62_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_55_cast <= SharedReg62_out;
SharedReg1073_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_56_cast <= SharedReg1073_out;
SharedReg1117_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1117_out;
SharedReg88_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_58_cast <= SharedReg88_out;
SharedReg1075_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_59_cast <= SharedReg1075_out;
SharedReg1119_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_60_cast <= SharedReg1119_out;
SharedReg1076_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_61_cast <= SharedReg1076_out;
SharedReg625_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_62_cast <= SharedReg625_out;
SharedReg266_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_63_cast <= SharedReg266_out;
SharedReg623_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_64_cast <= SharedReg623_out;
   MUX_Product31_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1079_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg624_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1087_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1088_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg235_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg235_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg909_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg88_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg618_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg618_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1093_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg89_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg913_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg619_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg954_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1106_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg88_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg617_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg617_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg88_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg932_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg89_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg621_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg95_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg92_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1061_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1062_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg623_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg937_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg265_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg623_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1137_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg97_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg914_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg75_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg270_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg272_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1067_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg275_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg100_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg628_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1097_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg629_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg944_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg944_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1083_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1101_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1070_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1071_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg906_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg62_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1073_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1117_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg88_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1075_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1119_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg607_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1076_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg625_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg266_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg623_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg236_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg247_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg105_out_to_MUX_Product31_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product31_2_impl_1_out);

   Delay1No77_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_2_impl_1_out,
                 Y => Delay1No77_out);

Delay1No78_out_to_Product31_3_impl_parent_implementedSystem_port_0_cast <= Delay1No78_out;
Delay1No79_out_to_Product31_3_impl_parent_implementedSystem_port_1_cast <= Delay1No79_out;
   Product31_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product31_3_impl_out,
                 X => Delay1No78_out_to_Product31_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No79_out_to_Product31_3_impl_parent_implementedSystem_port_1_cast);

SharedReg88_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg88_out;
SharedReg618_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg618_out;
SharedReg1074_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1074_out;
SharedReg115_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg115_out;
SharedReg641_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg641_out;
SharedReg267_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg267_out;
SharedReg1158_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1158_out;
SharedReg1077_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1077_out;
SharedReg1029_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1029_out;
SharedReg119_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg119_out;
SharedReg1159_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1159_out;
SharedReg1125_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1125_out;
SharedReg1081_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1081_out;
SharedReg1082_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1082_out;
SharedReg264_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg264_out;
SharedReg1084_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1084_out;
SharedReg1036_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1036_out;
SharedReg1037_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1037_out;
SharedReg1103_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1103_out;
SharedReg260_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg260_out;
SharedReg114_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg114_out;
SharedReg1089_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1089_out;
SharedReg1090_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1090_out;
SharedReg1145_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1145_out;
SharedReg1091_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1091_out;
SharedReg1132_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1132_out;
SharedReg1133_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1133_out;
SharedReg115_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg115_out;
SharedReg1094_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1094_out;
SharedReg1135_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1135_out;
SharedReg1105_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1105_out;
SharedReg110_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_32_cast <= SharedReg110_out;
SharedReg1046_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1046_out;
SharedReg1057_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1057_out;
SharedReg1170_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1170_out;
SharedReg1004_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1004_out;
SharedReg1166_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1166_out;
SharedReg1006_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1006_out;
SharedReg1171_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1171_out;
SharedReg1060_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1060_out;
SharedReg292_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_41_cast <= SharedReg292_out;
SharedReg290_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_42_cast <= SharedReg290_out;
SharedReg1115_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1115_out;
SharedReg1152_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1152_out;
SharedReg1063_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1063_out;
SharedReg1136_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1136_out;
SharedReg648_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_47_cast <= SharedReg648_out;
SharedReg1013_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1013_out;
SharedReg1120_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1120_out;
SharedReg1014_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1014_out;
SharedReg1015_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1015_out;
SharedReg296_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_52_cast <= SharedReg296_out;
SharedReg1017_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1017_out;
SharedReg1018_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1018_out;
SharedReg1047_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1047_out;
SharedReg124_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_56_cast <= SharedReg124_out;
SharedReg1049_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1049_out;
SharedReg1050_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1050_out;
SharedReg1051_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1051_out;
SharedReg269_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_60_cast <= SharedReg269_out;
SharedReg260_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_61_cast <= SharedReg260_out;
SharedReg640_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_62_cast <= SharedReg640_out;
SharedReg1156_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1156_out;
SharedReg1072_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1072_out;
   MUX_Product31_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg88_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg618_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1159_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1125_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1081_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1082_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg264_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1084_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1036_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1037_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1103_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg260_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1074_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg114_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1089_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1090_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1145_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1091_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1132_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1133_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg115_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1094_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1135_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg115_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1105_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg110_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1046_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1057_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1170_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1004_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1166_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1006_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1171_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1060_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg641_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg292_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg290_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1115_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1152_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1063_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1136_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg648_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1013_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1120_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1014_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg267_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1015_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg296_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1017_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1018_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1047_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg124_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1049_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1050_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1051_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg269_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1158_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg260_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg640_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1156_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1072_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1077_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1029_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg119_out_to_MUX_Product31_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product31_3_impl_0_out);

   Delay1No78_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_3_impl_0_out,
                 Y => Delay1No78_out);

SharedReg1073_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1073_out;
SharedReg1117_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1117_out;
SharedReg260_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg260_out;
SharedReg1075_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1075_out;
SharedReg1119_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1119_out;
SharedReg1076_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1076_out;
SharedReg939_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg939_out;
SharedReg119_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg119_out;
SharedReg937_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg937_out;
SharedReg1079_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1079_out;
SharedReg938_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg938_out;
SharedReg624_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg624_out;
SharedReg268_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg268_out;
SharedReg247_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg247_out;
SharedReg1083_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1083_out;
SharedReg920_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg920_out;
SharedReg262_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg262_out;
SharedReg100_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg100_out;
SharedReg130_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg130_out;
SharedReg1087_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1087_out;
SharedReg1088_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1088_out;
SharedReg261_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg261_out;
SharedReg261_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg261_out;
SharedReg934_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg934_out;
SharedReg114_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg114_out;
SharedReg641_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg641_out;
SharedReg641_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg641_out;
SharedReg1093_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1093_out;
SharedReg115_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_29_cast <= SharedReg115_out;
SharedReg642_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_30_cast <= SharedReg642_out;
SharedReg879_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_31_cast <= SharedReg879_out;
SharedReg1106_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_32_cast <= SharedReg1106_out;
SharedReg260_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_33_cast <= SharedReg260_out;
SharedReg640_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_34_cast <= SharedReg640_out;
SharedReg640_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_35_cast <= SharedReg640_out;
SharedReg114_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_36_cast <= SharedReg114_out;
SharedReg856_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_37_cast <= SharedReg856_out;
SharedReg115_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_38_cast <= SharedReg115_out;
SharedReg644_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_39_cast <= SharedReg644_out;
SharedReg118_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_40_cast <= SharedReg118_out;
SharedReg1061_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_41_cast <= SharedReg1061_out;
SharedReg1062_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_42_cast <= SharedReg1062_out;
SharedReg646_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_43_cast <= SharedReg646_out;
SharedReg861_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_44_cast <= SharedReg861_out;
SharedReg290_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_45_cast <= SharedReg290_out;
SharedReg646_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_46_cast <= SharedReg646_out;
SharedReg1137_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_47_cast <= SharedReg1137_out;
SharedReg123_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_48_cast <= SharedReg123_out;
SharedReg939_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_49_cast <= SharedReg939_out;
SharedReg295_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_50_cast <= SharedReg295_out;
SharedReg297_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_51_cast <= SharedReg297_out;
SharedReg1067_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_52_cast <= SharedReg1067_out;
SharedReg300_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_53_cast <= SharedReg300_out;
SharedReg125_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_54_cast <= SharedReg125_out;
SharedReg650_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_55_cast <= SharedReg650_out;
SharedReg1097_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_56_cast <= SharedReg1097_out;
SharedReg943_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_57_cast <= SharedReg943_out;
SharedReg869_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_58_cast <= SharedReg869_out;
SharedReg652_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_59_cast <= SharedReg652_out;
SharedReg1101_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_60_cast <= SharedReg1101_out;
SharedReg1070_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_61_cast <= SharedReg1070_out;
SharedReg1071_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_62_cast <= SharedReg1071_out;
SharedReg617_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_63_cast <= SharedReg617_out;
SharedReg234_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_64_cast <= SharedReg234_out;
   MUX_Product31_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1073_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1117_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg938_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg624_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg268_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg247_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1083_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg920_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg262_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg100_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg130_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1087_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg260_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1088_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg261_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg261_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg934_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg114_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg641_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg641_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1093_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg115_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg642_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1075_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg879_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1106_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg260_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg640_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg640_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg114_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg856_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg115_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg644_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg118_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1119_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1061_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1062_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg646_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg861_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg290_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg646_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1137_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg123_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg939_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg295_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1076_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg297_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1067_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg300_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg125_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg650_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1097_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg943_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg869_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg652_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1101_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg939_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1070_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1071_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg617_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg234_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg119_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg937_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1079_out_to_MUX_Product31_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product31_3_impl_1_out);

   Delay1No79_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_3_impl_1_out,
                 Y => Delay1No79_out);

Delay1No80_out_to_Product31_4_impl_parent_implementedSystem_port_0_cast <= Delay1No80_out;
Delay1No81_out_to_Product31_4_impl_parent_implementedSystem_port_1_cast <= Delay1No81_out;
   Product31_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product31_4_impl_out,
                 X => Delay1No80_out_to_Product31_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No81_out_to_Product31_4_impl_parent_implementedSystem_port_1_cast);

SharedReg149_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg149_out;
SharedReg1049_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1049_out;
SharedReg1050_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1050_out;
SharedReg1051_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1051_out;
SharedReg122_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg122_out;
SharedReg285_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg285_out;
SharedReg661_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg661_out;
SharedReg1156_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1156_out;
SharedReg1072_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1072_out;
SharedReg114_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg114_out;
SharedReg641_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg641_out;
SharedReg1074_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1074_out;
SharedReg140_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg140_out;
SharedReg662_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg662_out;
SharedReg292_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg292_out;
SharedReg1158_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1158_out;
SharedReg1077_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1077_out;
SharedReg1029_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1029_out;
SharedReg143_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg143_out;
SharedReg1159_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1159_out;
SharedReg1125_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1125_out;
SharedReg1081_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1081_out;
SharedReg1082_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1082_out;
SharedReg289_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg289_out;
SharedReg1084_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1084_out;
SharedReg1036_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1036_out;
SharedReg1037_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1037_out;
SharedReg1103_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1103_out;
SharedReg285_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_29_cast <= SharedReg285_out;
SharedReg139_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_30_cast <= SharedReg139_out;
SharedReg1089_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1089_out;
SharedReg1090_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1090_out;
SharedReg1145_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1145_out;
SharedReg1091_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1091_out;
SharedReg1132_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1132_out;
SharedReg1133_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1133_out;
SharedReg140_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_37_cast <= SharedReg140_out;
SharedReg1094_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1094_out;
SharedReg1135_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1135_out;
SharedReg1105_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1105_out;
SharedReg280_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_41_cast <= SharedReg280_out;
SharedReg1046_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1046_out;
SharedReg1057_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1057_out;
SharedReg1170_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1170_out;
SharedReg1004_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1004_out;
SharedReg1166_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1166_out;
SharedReg1006_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1006_out;
SharedReg1171_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1171_out;
SharedReg1060_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1060_out;
SharedReg316_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_50_cast <= SharedReg316_out;
SharedReg290_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_51_cast <= SharedReg290_out;
SharedReg1115_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1115_out;
SharedReg1152_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1152_out;
SharedReg1063_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1063_out;
SharedReg1136_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1136_out;
SharedReg669_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_56_cast <= SharedReg669_out;
SharedReg1013_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1013_out;
SharedReg1120_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1120_out;
SharedReg1014_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1014_out;
SharedReg1015_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1015_out;
SharedReg319_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_61_cast <= SharedReg319_out;
SharedReg1017_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1017_out;
SharedReg1018_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1018_out;
SharedReg1047_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1047_out;
   MUX_Product31_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg149_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1049_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg641_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1074_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg140_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg662_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg292_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1158_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1077_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1029_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg143_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1159_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1050_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1125_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1081_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1082_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg289_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1084_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1036_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1037_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1103_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg285_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg139_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1051_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1089_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1090_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1145_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1091_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1132_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1133_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg140_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1094_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1135_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1105_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg122_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg280_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1046_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1057_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1170_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1004_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1166_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1006_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1171_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1060_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg316_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg285_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg290_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1115_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1152_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1063_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1136_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg669_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1013_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1120_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1014_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1015_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg661_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg319_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1017_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1018_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1047_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1156_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1072_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg114_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product31_4_impl_0_out);

   Delay1No80_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_4_impl_0_out,
                 Y => Delay1No80_out);

SharedReg1097_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1097_out;
SharedReg867_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg867_out;
SharedReg698_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg698_out;
SharedReg675_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg675_out;
SharedReg1101_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1101_out;
SharedReg1070_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1070_out;
SharedReg1071_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1071_out;
SharedReg640_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg640_out;
SharedReg260_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg260_out;
SharedReg1073_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1073_out;
SharedReg1117_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1117_out;
SharedReg285_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg285_out;
SharedReg1075_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1075_out;
SharedReg1119_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1119_out;
SharedReg1076_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1076_out;
SharedReg863_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg863_out;
SharedReg143_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg143_out;
SharedReg861_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg861_out;
SharedReg1079_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1079_out;
SharedReg862_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg862_out;
SharedReg647_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg647_out;
SharedReg293_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg293_out;
SharedReg273_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg273_out;
SharedReg1083_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1083_out;
SharedReg945_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg945_out;
SharedReg287_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg287_out;
SharedReg125_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg125_out;
SharedReg305_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg305_out;
SharedReg1087_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_29_cast <= SharedReg1087_out;
SharedReg1088_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_30_cast <= SharedReg1088_out;
SharedReg286_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_31_cast <= SharedReg286_out;
SharedReg286_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_32_cast <= SharedReg286_out;
SharedReg858_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_33_cast <= SharedReg858_out;
SharedReg139_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_34_cast <= SharedReg139_out;
SharedReg662_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_35_cast <= SharedReg662_out;
SharedReg662_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_36_cast <= SharedReg662_out;
SharedReg1093_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_37_cast <= SharedReg1093_out;
SharedReg140_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_38_cast <= SharedReg140_out;
SharedReg663_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_39_cast <= SharedReg663_out;
SharedReg682_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_40_cast <= SharedReg682_out;
SharedReg1106_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_41_cast <= SharedReg1106_out;
SharedReg285_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_42_cast <= SharedReg285_out;
SharedReg661_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_43_cast <= SharedReg661_out;
SharedReg661_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_44_cast <= SharedReg661_out;
SharedReg285_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_45_cast <= SharedReg285_out;
SharedReg662_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_46_cast <= SharedReg662_out;
SharedReg115_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_47_cast <= SharedReg115_out;
SharedReg665_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_48_cast <= SharedReg665_out;
SharedReg142_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_49_cast <= SharedReg142_out;
SharedReg1061_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_50_cast <= SharedReg1061_out;
SharedReg1062_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_51_cast <= SharedReg1062_out;
SharedReg646_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_52_cast <= SharedReg646_out;
SharedReg667_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_53_cast <= SharedReg667_out;
SharedReg315_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_54_cast <= SharedReg315_out;
SharedReg667_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_55_cast <= SharedReg667_out;
SharedReg1137_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_56_cast <= SharedReg1137_out;
SharedReg295_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_57_cast <= SharedReg295_out;
SharedReg863_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_58_cast <= SharedReg863_out;
SharedReg318_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_59_cast <= SharedReg318_out;
SharedReg320_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_60_cast <= SharedReg320_out;
SharedReg1067_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_61_cast <= SharedReg1067_out;
SharedReg152_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_62_cast <= SharedReg152_out;
SharedReg150_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_63_cast <= SharedReg150_out;
SharedReg672_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_64_cast <= SharedReg672_out;
   MUX_Product31_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1097_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg867_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1117_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg285_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1075_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1119_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1076_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg863_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg143_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg861_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1079_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg862_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg698_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg647_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg293_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg273_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1083_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg945_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg287_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg125_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg305_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1087_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1088_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg675_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg286_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg286_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg858_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg139_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg662_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg662_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1093_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg140_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg663_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg682_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1101_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1106_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg285_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg661_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg661_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg285_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg662_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg115_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg665_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg142_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1061_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1070_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1062_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg646_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg667_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg315_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg667_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1137_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg295_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg863_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg318_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg320_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1071_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1067_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg152_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg150_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg672_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg640_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg260_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1073_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product31_4_impl_1_out);

   Delay1No81_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_4_impl_1_out,
                 Y => Delay1No81_out);

Delay1No82_out_to_Product31_5_impl_parent_implementedSystem_port_0_cast <= Delay1No82_out;
Delay1No83_out_to_Product31_5_impl_parent_implementedSystem_port_1_cast <= Delay1No83_out;
   Product31_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product31_5_impl_out,
                 X => Delay1No82_out_to_Product31_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No83_out_to_Product31_5_impl_parent_implementedSystem_port_1_cast);

SharedReg715_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg715_out;
SharedReg1013_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1013_out;
SharedReg1120_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1120_out;
SharedReg1014_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1014_out;
SharedReg1015_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1015_out;
SharedReg197_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg197_out;
SharedReg1017_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1017_out;
SharedReg1018_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1018_out;
SharedReg1047_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1047_out;
SharedReg320_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg320_out;
SharedReg1049_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1049_out;
SharedReg1050_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1050_out;
SharedReg1051_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1051_out;
SharedReg294_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_14_cast <= SharedReg294_out;
SharedReg310_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_15_cast <= SharedReg310_out;
SharedReg707_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_16_cast <= SharedReg707_out;
SharedReg1156_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1156_out;
SharedReg1072_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1072_out;
SharedReg139_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_19_cast <= SharedReg139_out;
SharedReg662_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_20_cast <= SharedReg662_out;
SharedReg1074_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1074_out;
SharedReg164_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_22_cast <= SharedReg164_out;
SharedReg708_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_23_cast <= SharedReg708_out;
SharedReg316_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_24_cast <= SharedReg316_out;
SharedReg1158_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1158_out;
SharedReg1077_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1077_out;
SharedReg1029_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1029_out;
SharedReg169_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_28_cast <= SharedReg169_out;
SharedReg1159_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1159_out;
SharedReg1125_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1125_out;
SharedReg1081_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1081_out;
SharedReg1082_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1082_out;
SharedReg314_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_33_cast <= SharedReg314_out;
SharedReg1084_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1084_out;
SharedReg1036_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1036_out;
SharedReg1037_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1037_out;
SharedReg1103_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1103_out;
SharedReg310_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_38_cast <= SharedReg310_out;
SharedReg163_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_39_cast <= SharedReg163_out;
SharedReg1089_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1089_out;
SharedReg1090_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1090_out;
SharedReg1145_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1145_out;
SharedReg1091_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1091_out;
SharedReg1132_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1132_out;
SharedReg1133_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1133_out;
SharedReg311_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_46_cast <= SharedReg311_out;
SharedReg1094_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1094_out;
SharedReg1135_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1135_out;
SharedReg1105_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1105_out;
SharedReg306_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_50_cast <= SharedReg306_out;
SharedReg1046_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1046_out;
SharedReg1057_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1057_out;
SharedReg1170_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1170_out;
SharedReg1004_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1004_out;
SharedReg1166_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1166_out;
SharedReg1006_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1006_out;
SharedReg1171_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1171_out;
SharedReg1060_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1060_out;
SharedReg193_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_59_cast <= SharedReg193_out;
SharedReg315_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_60_cast <= SharedReg315_out;
SharedReg1115_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1115_out;
SharedReg1152_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1152_out;
SharedReg1063_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1063_out;
SharedReg1136_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1136_out;
   MUX_Product31_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg715_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1013_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1049_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1050_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1051_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg294_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg310_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg707_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1156_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1072_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg139_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg662_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1120_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1074_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg164_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg708_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg316_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1158_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1077_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1029_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg169_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1159_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1125_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1014_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1081_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1082_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg314_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1084_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1036_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1037_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1103_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg310_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg163_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1089_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1015_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1090_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1145_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1091_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1132_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1133_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg311_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1094_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1135_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1105_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg306_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg197_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1046_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1057_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1170_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1004_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1166_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1006_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1171_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1060_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg193_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg315_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1017_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1115_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1152_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1063_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1136_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1018_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1047_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg320_out_to_MUX_Product31_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product31_5_impl_0_out);

   Delay1No82_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_5_impl_0_out,
                 Y => Delay1No82_out);

SharedReg1137_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1137_out;
SharedReg147_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg147_out;
SharedReg693_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg693_out;
SharedReg196_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg196_out;
SharedReg198_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg198_out;
SharedReg1067_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1067_out;
SharedReg323_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg323_out;
SharedReg175_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg175_out;
SharedReg696_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg696_out;
SharedReg1097_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1097_out;
SharedReg673_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg673_out;
SharedReg719_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg719_out;
SharedReg698_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg698_out;
SharedReg1101_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1101_out;
SharedReg1070_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1070_out;
SharedReg1071_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1071_out;
SharedReg661_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_17_cast <= SharedReg661_out;
SharedReg285_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_18_cast <= SharedReg285_out;
SharedReg1073_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1073_out;
SharedReg1117_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1117_out;
SharedReg310_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_21_cast <= SharedReg310_out;
SharedReg1075_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1075_out;
SharedReg1119_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_23_cast <= SharedReg1119_out;
SharedReg1076_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1076_out;
SharedReg693_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_25_cast <= SharedReg693_out;
SharedReg169_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_26_cast <= SharedReg169_out;
SharedReg691_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_27_cast <= SharedReg691_out;
SharedReg1079_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1079_out;
SharedReg692_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_29_cast <= SharedReg692_out;
SharedReg862_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_30_cast <= SharedReg862_out;
SharedReg317_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_31_cast <= SharedReg317_out;
SharedReg298_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_32_cast <= SharedReg298_out;
SharedReg1083_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_33_cast <= SharedReg1083_out;
SharedReg870_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_34_cast <= SharedReg870_out;
SharedReg141_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_35_cast <= SharedReg141_out;
SharedReg150_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_36_cast <= SharedReg150_out;
SharedReg327_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_37_cast <= SharedReg327_out;
SharedReg1087_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_38_cast <= SharedReg1087_out;
SharedReg1088_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_39_cast <= SharedReg1088_out;
SharedReg311_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_40_cast <= SharedReg311_out;
SharedReg311_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_41_cast <= SharedReg311_out;
SharedReg688_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_42_cast <= SharedReg688_out;
SharedReg163_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_43_cast <= SharedReg163_out;
SharedReg708_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_44_cast <= SharedReg708_out;
SharedReg708_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_45_cast <= SharedReg708_out;
SharedReg1093_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_46_cast <= SharedReg1093_out;
SharedReg140_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_47_cast <= SharedReg140_out;
SharedReg663_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_48_cast <= SharedReg663_out;
SharedReg726_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_49_cast <= SharedReg726_out;
SharedReg1106_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_50_cast <= SharedReg1106_out;
SharedReg310_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_51_cast <= SharedReg310_out;
SharedReg707_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_52_cast <= SharedReg707_out;
SharedReg707_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_53_cast <= SharedReg707_out;
SharedReg310_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_54_cast <= SharedReg310_out;
SharedReg708_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_55_cast <= SharedReg708_out;
SharedReg140_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_56_cast <= SharedReg140_out;
SharedReg711_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_57_cast <= SharedReg711_out;
SharedReg168_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_58_cast <= SharedReg168_out;
SharedReg1061_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_59_cast <= SharedReg1061_out;
SharedReg1062_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_60_cast <= SharedReg1062_out;
SharedReg667_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_61_cast <= SharedReg667_out;
SharedReg691_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_62_cast <= SharedReg691_out;
SharedReg191_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_63_cast <= SharedReg191_out;
SharedReg713_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_64_cast <= SharedReg713_out;
   MUX_Product31_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1137_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg147_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg673_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg719_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg698_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1101_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1070_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1071_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg661_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg285_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1073_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1117_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg693_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg310_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1075_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1119_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1076_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg693_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg169_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg691_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1079_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg692_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg862_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg196_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg317_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg298_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1083_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg870_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg141_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg150_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg327_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1087_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1088_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg311_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg198_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg311_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg688_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg163_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg708_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg708_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1093_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg140_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg663_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg726_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1106_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1067_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg310_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg707_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg707_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg310_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg708_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg140_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg711_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg168_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1061_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1062_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg323_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg667_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg691_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg191_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg713_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg175_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg696_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1097_out_to_MUX_Product31_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product31_5_impl_1_out);

   Delay1No83_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_5_impl_1_out,
                 Y => Delay1No83_out);

Delay1No84_out_to_Product31_6_impl_parent_implementedSystem_port_0_cast <= Delay1No84_out;
Delay1No85_out_to_Product31_6_impl_parent_implementedSystem_port_1_cast <= Delay1No85_out;
   Product31_6_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product31_6_impl_out,
                 X => Delay1No84_out_to_Product31_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No85_out_to_Product31_6_impl_parent_implementedSystem_port_1_cast);

SharedReg1166_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1166_out;
SharedReg1006_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1006_out;
SharedReg1171_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1171_out;
SharedReg1060_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1060_out;
SharedReg339_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg339_out;
SharedReg168_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg168_out;
SharedReg1115_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1115_out;
SharedReg1152_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1152_out;
SharedReg1063_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1063_out;
SharedReg1136_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1136_out;
SharedReg890_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg890_out;
SharedReg1013_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1013_out;
SharedReg1120_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1120_out;
SharedReg1014_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1014_out;
SharedReg1015_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1015_out;
SharedReg173_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_16_cast <= SharedReg173_out;
SharedReg1017_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1017_out;
SharedReg1018_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1018_out;
SharedReg1047_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1047_out;
SharedReg174_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_20_cast <= SharedReg174_out;
SharedReg1049_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1049_out;
SharedReg1050_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1050_out;
SharedReg1051_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1051_out;
SharedReg195_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_24_cast <= SharedReg195_out;
SharedReg186_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_25_cast <= SharedReg186_out;
SharedReg882_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_26_cast <= SharedReg882_out;
SharedReg1156_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1156_out;
SharedReg1072_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1072_out;
SharedReg332_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_29_cast <= SharedReg332_out;
SharedReg984_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_30_cast <= SharedReg984_out;
SharedReg1074_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1074_out;
SharedReg333_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_32_cast <= SharedReg333_out;
SharedReg708_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_33_cast <= SharedReg708_out;
SharedReg170_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_34_cast <= SharedReg170_out;
SharedReg1158_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1158_out;
SharedReg1077_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1077_out;
SharedReg1029_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1029_out;
SharedReg192_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_38_cast <= SharedReg192_out;
SharedReg1159_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1159_out;
SharedReg1125_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1125_out;
SharedReg1081_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1081_out;
SharedReg1082_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1082_out;
SharedReg190_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_43_cast <= SharedReg190_out;
SharedReg1084_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1084_out;
SharedReg1036_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1036_out;
SharedReg1037_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1037_out;
SharedReg1103_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1103_out;
SharedReg186_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_48_cast <= SharedReg186_out;
SharedReg332_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_49_cast <= SharedReg332_out;
SharedReg1089_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1089_out;
SharedReg1090_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1090_out;
SharedReg1145_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1145_out;
SharedReg1091_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1091_out;
SharedReg1132_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1132_out;
SharedReg1133_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1133_out;
SharedReg164_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_56_cast <= SharedReg164_out;
SharedReg1094_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1094_out;
SharedReg1135_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1135_out;
SharedReg1105_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1105_out;
SharedReg205_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_60_cast <= SharedReg205_out;
SharedReg1046_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1046_out;
SharedReg1057_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1057_out;
SharedReg1170_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1170_out;
SharedReg1004_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1004_out;
   MUX_Product31_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1166_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1006_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg890_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1013_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1120_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1014_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1015_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg173_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1017_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1018_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1047_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg174_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1171_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1049_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1050_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1051_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg195_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg186_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg882_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1156_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1072_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg332_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg984_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1060_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1074_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg333_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg708_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg170_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1158_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1077_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1029_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg192_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1159_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1125_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg339_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1081_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1082_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg190_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1084_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1036_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1037_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1103_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg186_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg332_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1089_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg168_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1090_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1145_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1091_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1132_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1133_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg164_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1094_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1135_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1105_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg205_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1115_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1046_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1057_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1170_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1004_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1152_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1063_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1136_out_to_MUX_Product31_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product31_6_impl_0_out);

   Delay1No84_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_6_impl_0_out,
                 Y => Delay1No84_out);

SharedReg708_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg708_out;
SharedReg311_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg311_out;
SharedReg711_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg711_out;
SharedReg168_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg168_out;
SharedReg1061_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1061_out;
SharedReg1062_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1062_out;
SharedReg691_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg691_out;
SharedReg989_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg989_out;
SharedReg337_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg337_out;
SharedReg713_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg713_out;
SharedReg1137_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1137_out;
SharedReg196_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg196_out;
SharedReg715_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_13_cast <= SharedReg715_out;
SharedReg341_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_14_cast <= SharedReg341_out;
SharedReg342_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_15_cast <= SharedReg342_out;
SharedReg1067_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1067_out;
SharedReg343_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_17_cast <= SharedReg343_out;
SharedReg321_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_18_cast <= SharedReg321_out;
SharedReg717_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_19_cast <= SharedReg717_out;
SharedReg1097_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1097_out;
SharedReg697_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_21_cast <= SharedReg697_out;
SharedReg895_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_22_cast <= SharedReg895_out;
SharedReg719_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_23_cast <= SharedReg719_out;
SharedReg1101_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1101_out;
SharedReg1070_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1070_out;
SharedReg1071_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1071_out;
SharedReg685_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_27_cast <= SharedReg685_out;
SharedReg310_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_28_cast <= SharedReg310_out;
SharedReg1073_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_29_cast <= SharedReg1073_out;
SharedReg1117_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_30_cast <= SharedReg1117_out;
SharedReg186_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_31_cast <= SharedReg186_out;
SharedReg1075_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_32_cast <= SharedReg1075_out;
SharedReg1119_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_33_cast <= SharedReg1119_out;
SharedReg1076_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_34_cast <= SharedReg1076_out;
SharedReg715_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_35_cast <= SharedReg715_out;
SharedReg338_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_36_cast <= SharedReg338_out;
SharedReg888_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_37_cast <= SharedReg888_out;
SharedReg1079_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_38_cast <= SharedReg1079_out;
SharedReg692_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_39_cast <= SharedReg692_out;
SharedReg889_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_40_cast <= SharedReg889_out;
SharedReg194_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_41_cast <= SharedReg194_out;
SharedReg199_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_42_cast <= SharedReg199_out;
SharedReg1083_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_43_cast <= SharedReg1083_out;
SharedReg896_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_44_cast <= SharedReg896_out;
SharedReg188_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_45_cast <= SharedReg188_out;
SharedReg175_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_46_cast <= SharedReg175_out;
SharedReg178_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_47_cast <= SharedReg178_out;
SharedReg1087_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_48_cast <= SharedReg1087_out;
SharedReg1088_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_49_cast <= SharedReg1088_out;
SharedReg187_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_50_cast <= SharedReg187_out;
SharedReg187_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_51_cast <= SharedReg187_out;
SharedReg885_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_52_cast <= SharedReg885_out;
SharedReg332_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_53_cast <= SharedReg332_out;
SharedReg984_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_54_cast <= SharedReg984_out;
SharedReg883_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_55_cast <= SharedReg883_out;
SharedReg1093_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_56_cast <= SharedReg1093_out;
SharedReg164_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_57_cast <= SharedReg164_out;
SharedReg709_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_58_cast <= SharedReg709_out;
SharedReg1000_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_59_cast <= SharedReg1000_out;
SharedReg1106_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_60_cast <= SharedReg1106_out;
SharedReg186_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_61_cast <= SharedReg186_out;
SharedReg882_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_62_cast <= SharedReg882_out;
SharedReg707_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_63_cast <= SharedReg707_out;
SharedReg310_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_64_cast <= SharedReg310_out;
   MUX_Product31_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg708_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg311_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1137_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg196_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg715_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg341_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg342_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1067_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg343_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg321_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg717_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1097_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg711_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg697_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg895_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg719_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1101_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1070_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1071_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg685_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg310_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1073_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1117_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg168_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg186_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1075_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1119_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1076_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg715_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg338_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg888_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1079_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg692_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg889_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1061_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg194_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg199_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1083_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg896_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg188_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg175_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg178_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1087_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1088_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg187_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1062_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg187_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg885_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg332_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg984_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg883_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1093_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg164_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg709_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1000_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1106_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg691_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg186_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg882_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg707_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg310_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg989_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg337_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg713_out_to_MUX_Product31_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product31_6_impl_1_out);

   Delay1No85_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_6_impl_1_out,
                 Y => Delay1No85_out);

Delay1No86_out_to_Subtract2_0_impl_parent_implementedSystem_port_0_cast <= Delay1No86_out;
Delay1No87_out_to_Subtract2_0_impl_parent_implementedSystem_port_1_cast <= Delay1No87_out;
   Subtract2_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_0_impl_out,
                 X => Delay1No86_out_to_Subtract2_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No87_out_to_Subtract2_0_impl_parent_implementedSystem_port_1_cast);

SharedReg350_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg350_out;
SharedReg_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg_out;
SharedReg2_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg2_out;
SharedReg14_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg14_out;
SharedReg4_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg7_out;
SharedReg10_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg10_out;
SharedReg9_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg9_out;
SharedReg8_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg8_out;
SharedReg358_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg358_out;
SharedReg355_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg355_out;
SharedReg52_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg52_out;
SharedReg582_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg582_out;
SharedReg467_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg467_out;
SharedReg455_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg455_out;
SharedReg737_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg737_out;
SharedReg743_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg743_out;
SharedReg356_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg356_out;
SharedReg730_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg730_out;
SharedReg350_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg350_out;
SharedReg729_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg729_out;
SharedReg959_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg959_out;
SharedReg38_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg38_out;
SharedReg351_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg351_out;
SharedReg211_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg211_out;
SharedReg350_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg350_out;
SharedReg356_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg356_out;
SharedReg963_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg963_out;
SharedReg458_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_29_cast <= SharedReg458_out;
SharedReg455_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_30_cast <= SharedReg455_out;
SharedReg567_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_31_cast <= SharedReg567_out;
SharedReg350_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_32_cast <= SharedReg350_out;
SharedReg961_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_33_cast <= SharedReg961_out;
SharedReg208_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_34_cast <= SharedReg208_out;
SharedReg48_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_35_cast <= SharedReg48_out;
SharedReg569_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_36_cast <= SharedReg569_out;
SharedReg53_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_37_cast <= SharedReg53_out;
SharedReg354_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_38_cast <= SharedReg354_out;
SharedReg459_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_39_cast <= SharedReg459_out;
SharedReg458_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_40_cast <= SharedReg458_out;
SharedReg365_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_41_cast <= SharedReg365_out;
SharedReg351_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_42_cast <= SharedReg351_out;
SharedReg730_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_43_cast <= SharedReg730_out;
SharedReg583_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_44_cast <= SharedReg583_out;
SharedReg351_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_45_cast <= SharedReg351_out;
SharedReg730_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_46_cast <= SharedReg730_out;
SharedReg39_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_47_cast <= SharedReg39_out;
SharedReg350_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_48_cast <= SharedReg350_out;
SharedReg213_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_49_cast <= SharedReg213_out;
SharedReg350_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_50_cast <= SharedReg350_out;
SharedReg352_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_51_cast <= SharedReg352_out;
SharedReg455_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_52_cast <= SharedReg455_out;
SharedReg573_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_53_cast <= SharedReg573_out;
SharedReg352_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_54_cast <= SharedReg352_out;
SharedReg350_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_55_cast <= SharedReg350_out;
SharedReg352_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_56_cast <= SharedReg352_out;
SharedReg573_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_57_cast <= SharedReg573_out;
SharedReg215_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_58_cast <= SharedReg215_out;
SharedReg217_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_59_cast <= SharedReg217_out;
SharedReg576_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_60_cast <= SharedReg576_out;
SharedReg735_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_61_cast <= SharedReg735_out;
SharedReg355_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_62_cast <= SharedReg355_out;
SharedReg350_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_63_cast <= SharedReg350_out;
SharedReg350_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_64_cast <= SharedReg350_out;
   MUX_Subtract2_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg350_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg355_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg52_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg582_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg467_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg455_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg737_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg743_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg356_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg730_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg350_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg2_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg729_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg959_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg38_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg351_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg211_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg350_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg356_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg963_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg458_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg455_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg14_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg567_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg350_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg961_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg208_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg48_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg569_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg53_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg354_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg459_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg458_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg4_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg365_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg351_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg730_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg583_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg351_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg730_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg39_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg350_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg213_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg350_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg7_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg352_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg455_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg573_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg352_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg350_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg352_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg573_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg215_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg217_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg576_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg10_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg735_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg355_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg350_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg350_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg9_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg8_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg358_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract2_0_impl_0_out);

   Delay1No86_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_0_impl_0_out,
                 Y => Delay1No86_out);

SharedReg733_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg733_out;
SharedReg18_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg20_out;
SharedReg32_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg32_out;
SharedReg22_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg25_out;
SharedReg28_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg28_out;
SharedReg27_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg27_out;
SharedReg26_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg26_out;
SharedReg357_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg357_out;
SharedReg460_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg460_out;
SharedReg51_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg51_out;
SharedReg581_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg581_out;
SharedReg362_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg362_out;
SharedReg731_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg731_out;
Delay44No_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_16_cast <= Delay44No_out;
SharedReg462_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg462_out;
SharedReg455_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg455_out;
SharedReg350_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg350_out;
SharedReg732_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg732_out;
SharedReg358_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg358_out;
SharedReg591_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg591_out;
SharedReg232_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg232_out;
SharedReg455_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg455_out;
SharedReg61_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg61_out;
SharedReg351_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg351_out;
SharedReg350_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg350_out;
Delay78No_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_28_cast <= Delay78No_out;
SharedReg455_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_29_cast <= SharedReg455_out;
SharedReg731_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_30_cast <= SharedReg731_out;
SharedReg572_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_31_cast <= SharedReg572_out;
SharedReg360_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_32_cast <= SharedReg360_out;
SharedReg571_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_33_cast <= SharedReg571_out;
SharedReg210_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_34_cast <= SharedReg210_out;
SharedReg36_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_35_cast <= SharedReg36_out;
SharedReg961_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_36_cast <= SharedReg961_out;
SharedReg208_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_37_cast <= SharedReg208_out;
SharedReg745_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_38_cast <= SharedReg745_out;
SharedReg736_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_39_cast <= SharedReg736_out;
SharedReg734_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_40_cast <= SharedReg734_out;
SharedReg375_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_41_cast <= SharedReg375_out;
SharedReg455_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_42_cast <= SharedReg455_out;
SharedReg455_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_43_cast <= SharedReg455_out;
SharedReg958_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_44_cast <= SharedReg958_out;
SharedReg455_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_45_cast <= SharedReg455_out;
SharedReg455_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_46_cast <= SharedReg455_out;
SharedReg228_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_47_cast <= SharedReg228_out;
SharedReg456_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_48_cast <= SharedReg456_out;
SharedReg59_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_49_cast <= SharedReg59_out;
SharedReg730_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_50_cast <= SharedReg730_out;
SharedReg455_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_51_cast <= SharedReg455_out;
SharedReg738_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_52_cast <= SharedReg738_out;
SharedReg567_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_53_cast <= SharedReg567_out;
SharedReg732_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_54_cast <= SharedReg732_out;
SharedReg465_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_55_cast <= SharedReg465_out;
SharedReg455_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_56_cast <= SharedReg455_out;
SharedReg567_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_57_cast <= SharedReg567_out;
SharedReg209_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_58_cast <= SharedReg209_out;
SharedReg208_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_59_cast <= SharedReg208_out;
SharedReg568_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_60_cast <= SharedReg568_out;
SharedReg733_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_61_cast <= SharedReg733_out;
SharedReg468_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_62_cast <= SharedReg468_out;
SharedReg457_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_63_cast <= SharedReg457_out;
SharedReg457_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_64_cast <= SharedReg457_out;
   MUX_Subtract2_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg733_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg18_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg460_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg51_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg581_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg362_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg731_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => Delay44No_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg462_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg455_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg350_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg732_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg20_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg358_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg591_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg232_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg455_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg61_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg351_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg350_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => Delay78No_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg455_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg731_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg32_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg572_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg360_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg571_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg210_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg36_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg961_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg208_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg745_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg736_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg734_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg22_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg375_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg455_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg455_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg958_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg455_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg455_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg228_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg456_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg59_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg730_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg25_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg455_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg738_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg567_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg732_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg465_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg455_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg567_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg209_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg208_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg568_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg28_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg733_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg468_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg457_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg457_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg27_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg26_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg357_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract2_0_impl_1_out);

   Delay1No87_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_0_impl_1_out,
                 Y => Delay1No87_out);

Delay1No88_out_to_Subtract2_1_impl_parent_implementedSystem_port_0_cast <= Delay1No88_out;
Delay1No89_out_to_Subtract2_1_impl_parent_implementedSystem_port_1_cast <= Delay1No89_out;
   Subtract2_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_1_impl_out,
                 X => Delay1No88_out_to_Subtract2_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No89_out_to_Subtract2_1_impl_parent_implementedSystem_port_1_cast);

SharedReg367_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg367_out;
SharedReg963_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg963_out;
SharedReg69_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg69_out;
SharedReg243_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg243_out;
SharedReg602_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg602_out;
SharedReg753_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg753_out;
SharedReg370_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg370_out;
SharedReg365_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg365_out;
SharedReg365_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg365_out;
SharedReg365_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg365_out;
SharedReg_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg_out;
SharedReg2_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg2_out;
SharedReg14_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg14_out;
SharedReg4_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg7_out;
SharedReg10_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg10_out;
SharedReg9_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg9_out;
SharedReg13_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg13_out;
SharedReg373_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg373_out;
SharedReg370_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg370_out;
SharedReg224_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg224_out;
SharedReg973_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg973_out;
SharedReg483_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg483_out;
SharedReg471_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg471_out;
SharedReg755_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg755_out;
SharedReg761_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg761_out;
SharedReg371_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg371_out;
SharedReg748_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg748_out;
SharedReg365_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_29_cast <= SharedReg365_out;
SharedReg747_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_30_cast <= SharedReg747_out;
SharedReg908_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_31_cast <= SharedReg908_out;
SharedReg64_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_32_cast <= SharedReg64_out;
SharedReg366_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_33_cast <= SharedReg366_out;
SharedReg237_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_34_cast <= SharedReg237_out;
SharedReg365_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_35_cast <= SharedReg365_out;
SharedReg371_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_36_cast <= SharedReg371_out;
SharedReg912_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_37_cast <= SharedReg912_out;
SharedReg474_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_38_cast <= SharedReg474_out;
SharedReg471_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_39_cast <= SharedReg471_out;
SharedReg234_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_40_cast <= SharedReg234_out;
SharedReg90_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_41_cast <= SharedReg90_out;
SharedReg246_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_42_cast <= SharedReg246_out;
SharedReg234_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_43_cast <= SharedReg234_out;
SharedReg74_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_44_cast <= SharedReg74_out;
SharedReg595_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_45_cast <= SharedReg595_out;
SharedReg78_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_46_cast <= SharedReg78_out;
SharedReg369_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_47_cast <= SharedReg369_out;
SharedReg475_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_48_cast <= SharedReg475_out;
SharedReg474_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_49_cast <= SharedReg474_out;
SharedReg380_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_50_cast <= SharedReg380_out;
SharedReg621_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_51_cast <= SharedReg621_out;
SharedReg748_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_52_cast <= SharedReg748_out;
SharedReg609_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_53_cast <= SharedReg609_out;
SharedReg366_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_54_cast <= SharedReg366_out;
SharedReg595_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_55_cast <= SharedReg595_out;
SharedReg909_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_56_cast <= SharedReg909_out;
SharedReg478_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_57_cast <= SharedReg478_out;
SharedReg597_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_58_cast <= SharedReg597_out;
SharedReg67_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_59_cast <= SharedReg67_out;
SharedReg381_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_60_cast <= SharedReg381_out;
SharedReg213_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_61_cast <= SharedReg213_out;
SharedReg239_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_62_cast <= SharedReg239_out;
SharedReg599_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_63_cast <= SharedReg599_out;
SharedReg766_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_64_cast <= SharedReg766_out;
   MUX_Subtract2_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg367_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg963_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg2_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg14_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg4_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg7_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg10_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg9_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg13_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg373_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg370_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg69_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg224_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg973_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg483_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg471_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg755_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg761_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg371_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg748_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg365_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg747_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg243_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg908_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg64_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg366_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg237_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg365_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg371_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg912_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg474_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg471_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg234_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg602_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg90_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg246_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg234_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg74_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg595_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg78_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg369_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg475_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg474_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg380_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg753_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg621_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg748_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg609_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg366_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg595_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg909_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg478_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg597_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg67_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg381_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg370_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg213_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg239_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg599_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg766_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg365_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg365_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg365_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract2_1_impl_0_out);

   Delay1No88_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_1_impl_0_out,
                 Y => Delay1No88_out);

SharedReg471_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg471_out;
SharedReg957_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg957_out;
SharedReg63_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg63_out;
SharedReg62_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg62_out;
SharedReg958_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg958_out;
SharedReg751_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg751_out;
SharedReg484_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg484_out;
SharedReg473_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg473_out;
SharedReg473_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg473_out;
SharedReg751_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg751_out;
SharedReg18_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg20_out;
SharedReg32_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg32_out;
SharedReg22_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg25_out;
SharedReg28_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg28_out;
SharedReg27_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg27_out;
SharedReg31_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg31_out;
SharedReg372_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg372_out;
SharedReg476_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg476_out;
SharedReg77_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg77_out;
SharedReg608_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg608_out;
SharedReg377_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg377_out;
SharedReg749_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg749_out;
Delay44No1_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_25_cast <= Delay44No1_out;
SharedReg478_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg478_out;
SharedReg471_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg471_out;
SharedReg365_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg365_out;
SharedReg750_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_29_cast <= SharedReg750_out;
SharedReg373_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_30_cast <= SharedReg373_out;
SharedReg615_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_31_cast <= SharedReg615_out;
SharedReg257_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_32_cast <= SharedReg257_out;
SharedReg471_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_33_cast <= SharedReg471_out;
SharedReg87_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_34_cast <= SharedReg87_out;
SharedReg366_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_35_cast <= SharedReg366_out;
SharedReg365_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_36_cast <= SharedReg365_out;
Delay78No1_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_37_cast <= Delay78No1_out;
SharedReg471_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_38_cast <= SharedReg471_out;
SharedReg749_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_39_cast <= SharedReg749_out;
SharedReg240_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_40_cast <= SharedReg240_out;
SharedReg282_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_41_cast <= SharedReg282_out;
SharedReg62_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_42_cast <= SharedReg62_out;
SharedReg236_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_43_cast <= SharedReg236_out;
SharedReg62_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_44_cast <= SharedReg62_out;
SharedReg910_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_45_cast <= SharedReg910_out;
SharedReg208_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_46_cast <= SharedReg208_out;
SharedReg763_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_47_cast <= SharedReg763_out;
SharedReg754_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_48_cast <= SharedReg754_out;
SharedReg752_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_49_cast <= SharedReg752_out;
SharedReg390_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_50_cast <= SharedReg390_out;
SharedReg910_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_51_cast <= SharedReg910_out;
SharedReg471_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_52_cast <= SharedReg471_out;
SharedReg907_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_53_cast <= SharedReg907_out;
SharedReg471_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_54_cast <= SharedReg471_out;
SharedReg612_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_55_cast <= SharedReg612_out;
SharedReg613_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_56_cast <= SharedReg613_out;
SharedReg747_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_57_cast <= SharedReg747_out;
SharedReg928_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_58_cast <= SharedReg928_out;
SharedReg256_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_59_cast <= SharedReg256_out;
SharedReg487_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_60_cast <= SharedReg487_out;
SharedReg62_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_61_cast <= SharedReg62_out;
SharedReg62_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_62_cast <= SharedReg62_out;
SharedReg594_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_63_cast <= SharedReg594_out;
SharedReg487_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_64_cast <= SharedReg487_out;
   MUX_Subtract2_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg471_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg957_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg18_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg20_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg32_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg22_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg25_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg28_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg27_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg31_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg372_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg476_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg63_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg77_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg608_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg377_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg749_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => Delay44No1_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg478_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg471_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg365_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg750_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg373_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg62_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg615_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg257_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg471_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg87_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg366_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg365_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => Delay78No1_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg471_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg749_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg240_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg958_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg282_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg62_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg236_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg62_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg910_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg208_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg763_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg754_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg752_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg390_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg751_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg910_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg471_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg907_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg471_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg612_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg613_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg747_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg928_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg256_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg487_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg484_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg62_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg62_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg594_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg487_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg473_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg473_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg751_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract2_1_impl_1_out);

   Delay1No89_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_1_impl_1_out,
                 Y => Delay1No89_out);

Delay1No90_out_to_Subtract2_2_impl_parent_implementedSystem_port_0_cast <= Delay1No90_out;
Delay1No91_out_to_Subtract2_2_impl_parent_implementedSystem_port_1_cast <= Delay1No91_out;
   Subtract2_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_2_impl_out,
                 X => Delay1No90_out_to_Subtract2_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No91_out_to_Subtract2_2_impl_parent_implementedSystem_port_1_cast);

SharedReg620_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg620_out;
SharedReg494_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg494_out;
SharedReg910_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg910_out;
SharedReg239_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg239_out;
SharedReg396_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg396_out;
SharedReg67_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg67_out;
SharedReg92_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg92_out;
SharedReg912_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg912_out;
SharedReg784_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg784_out;
SharedReg382_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg382_out;
SharedReg599_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg599_out;
SharedReg241_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg241_out;
SharedReg96_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg96_out;
SharedReg916_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg916_out;
SharedReg771_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg771_out;
SharedReg385_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg385_out;
SharedReg380_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg380_out;
SharedReg395_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg395_out;
SharedReg380_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg380_out;
SharedReg_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg_out;
SharedReg2_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg2_out;
SharedReg14_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg14_out;
SharedReg4_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg7_out;
SharedReg10_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg10_out;
SharedReg9_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg9_out;
SharedReg13_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg13_out;
SharedReg388_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg388_out;
SharedReg385_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_29_cast <= SharedReg385_out;
SharedReg250_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_30_cast <= SharedReg250_out;
SharedReg921_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_31_cast <= SharedReg921_out;
SharedReg499_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_32_cast <= SharedReg499_out;
SharedReg487_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_33_cast <= SharedReg487_out;
SharedReg773_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_34_cast <= SharedReg773_out;
SharedReg779_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_35_cast <= SharedReg779_out;
SharedReg386_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_36_cast <= SharedReg386_out;
SharedReg766_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_37_cast <= SharedReg766_out;
SharedReg380_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_38_cast <= SharedReg380_out;
SharedReg765_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_39_cast <= SharedReg765_out;
SharedReg262_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_40_cast <= SharedReg262_out;
SharedReg515_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_41_cast <= SharedReg515_out;
SharedReg765_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_42_cast <= SharedReg765_out;
SharedReg263_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_43_cast <= SharedReg263_out;
SharedReg380_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_44_cast <= SharedReg380_out;
SharedReg386_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_45_cast <= SharedReg386_out;
SharedReg937_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_46_cast <= SharedReg937_out;
SharedReg490_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_47_cast <= SharedReg490_out;
SharedReg487_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_48_cast <= SharedReg487_out;
SharedReg260_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_49_cast <= SharedReg260_out;
SharedReg116_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_50_cast <= SharedReg116_out;
SharedReg396_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_51_cast <= SharedReg396_out;
SharedReg260_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_52_cast <= SharedReg260_out;
SharedReg99_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_53_cast <= SharedReg99_out;
SharedReg619_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_54_cast <= SharedReg619_out;
SharedReg630_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_55_cast <= SharedReg630_out;
SharedReg493_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_56_cast <= SharedReg493_out;
SharedReg383_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_57_cast <= SharedReg383_out;
SharedReg640_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_58_cast <= SharedReg640_out;
SharedReg866_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_59_cast <= SharedReg866_out;
SharedReg297_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_60_cast <= SharedReg297_out;
SharedReg104_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_61_cast <= SharedReg104_out;
SharedReg907_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_62_cast <= SharedReg907_out;
SharedReg90_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_63_cast <= SharedReg90_out;
SharedReg277_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_64_cast <= SharedReg277_out;
   MUX_Subtract2_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg620_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg494_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg599_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg241_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg96_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg916_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg771_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg385_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg380_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg395_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg380_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg910_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg2_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg14_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg4_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg7_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg10_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg9_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg13_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg388_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg385_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg250_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg239_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg921_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg499_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg487_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg773_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg779_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg386_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg766_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg380_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg765_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg262_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg396_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg515_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg765_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg263_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg380_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg386_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg937_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg490_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg487_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg260_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg116_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg67_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg396_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg260_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg99_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg619_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg630_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg493_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg383_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg640_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg866_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg297_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg92_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg104_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg907_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg90_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg277_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg912_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg784_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg382_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract2_2_impl_0_out);

   Delay1No90_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_2_impl_0_out,
                 Y => Delay1No90_out);

SharedReg927_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg927_out;
SharedReg765_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg765_out;
SharedReg954_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg954_out;
SharedReg281_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg281_out;
SharedReg503_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg503_out;
SharedReg88_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg88_out;
SharedReg88_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg88_out;
SharedReg618_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg618_out;
SharedReg503_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg503_out;
SharedReg487_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg487_out;
SharedReg906_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg906_out;
SharedReg89_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg89_out;
SharedReg88_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg88_out;
SharedReg907_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg907_out;
SharedReg769_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg769_out;
SharedReg500_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg500_out;
SharedReg489_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg489_out;
SharedReg513_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg513_out;
SharedReg769_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg769_out;
SharedReg18_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg20_out;
SharedReg32_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg32_out;
SharedReg22_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg25_out;
SharedReg28_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg28_out;
SharedReg27_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg27_out;
SharedReg31_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg31_out;
SharedReg387_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg387_out;
SharedReg492_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_29_cast <= SharedReg492_out;
SharedReg102_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_30_cast <= SharedReg102_out;
SharedReg632_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_31_cast <= SharedReg632_out;
SharedReg392_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_32_cast <= SharedReg392_out;
SharedReg767_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_33_cast <= SharedReg767_out;
Delay44No2_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_34_cast <= Delay44No2_out;
SharedReg494_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_35_cast <= SharedReg494_out;
SharedReg487_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_36_cast <= SharedReg487_out;
SharedReg380_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_37_cast <= SharedReg380_out;
SharedReg768_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_38_cast <= SharedReg768_out;
SharedReg388_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_39_cast <= SharedReg388_out;
SharedReg113_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_40_cast <= SharedReg113_out;
SharedReg407_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_41_cast <= SharedReg407_out;
SharedReg775_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_42_cast <= SharedReg775_out;
SharedReg258_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_43_cast <= SharedReg258_out;
SharedReg381_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_44_cast <= SharedReg381_out;
SharedReg380_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_45_cast <= SharedReg380_out;
Delay78No2_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_46_cast <= Delay78No2_out;
SharedReg487_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_47_cast <= SharedReg487_out;
SharedReg767_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_48_cast <= SharedReg767_out;
SharedReg266_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_49_cast <= SharedReg266_out;
SharedReg307_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_50_cast <= SharedReg307_out;
SharedReg503_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_51_cast <= SharedReg503_out;
SharedReg262_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_52_cast <= SharedReg262_out;
SharedReg88_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_53_cast <= SharedReg88_out;
SharedReg935_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_54_cast <= SharedReg935_out;
SharedReg593_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_55_cast <= SharedReg593_out;
SharedReg498_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_56_cast <= SharedReg498_out;
SharedReg492_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_57_cast <= SharedReg492_out;
SharedReg645_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_58_cast <= SharedReg645_out;
SharedReg640_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_59_cast <= SharedReg640_out;
SharedReg260_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_60_cast <= SharedReg260_out;
SharedReg234_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_61_cast <= SharedReg234_out;
SharedReg637_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_62_cast <= SharedReg637_out;
SharedReg111_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_63_cast <= SharedReg111_out;
SharedReg88_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_64_cast <= SharedReg88_out;
   MUX_Subtract2_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg927_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg765_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg906_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg89_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg88_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg907_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg769_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg500_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg489_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg513_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg769_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg18_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg954_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg20_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg32_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg22_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg25_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg28_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg27_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg31_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg387_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg492_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg102_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg281_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg632_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg392_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg767_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => Delay44No2_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg494_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg487_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg380_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg768_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg388_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg113_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg503_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg407_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg775_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg258_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg381_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg380_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => Delay78No2_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg487_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg767_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg266_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg307_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg88_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg503_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg262_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg88_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg935_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg593_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg498_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg492_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg645_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg640_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg260_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg88_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg234_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg637_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg111_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg88_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg618_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg503_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg487_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract2_2_impl_1_out);

   Delay1No91_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_2_impl_1_out,
                 Y => Delay1No91_out);

Delay1No92_out_to_Subtract2_3_impl_parent_implementedSystem_port_0_cast <= Delay1No92_out;
Delay1No93_out_to_Subtract2_3_impl_parent_implementedSystem_port_1_cast <= Delay1No93_out;
   Subtract2_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_3_impl_out,
                 X => Delay1No92_out_to_Subtract2_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No93_out_to_Subtract2_3_impl_parent_implementedSystem_port_1_cast);

SharedReg509_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg509_out;
SharedReg398_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg398_out;
SharedReg855_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg855_out;
SharedReg696_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg696_out;
SharedReg320_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg320_out;
SharedReg129_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg129_out;
SharedReg932_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg932_out;
SharedReg116_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg116_out;
SharedReg128_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg128_out;
SharedReg643_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg643_out;
SharedReg510_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg510_out;
SharedReg935_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg935_out;
SharedReg265_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg265_out;
SharedReg411_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg411_out;
SharedReg92_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg92_out;
SharedReg118_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg118_out;
SharedReg937_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg937_out;
SharedReg857_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg857_out;
SharedReg397_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg397_out;
SharedReg623_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg623_out;
SharedReg267_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg267_out;
SharedReg122_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg122_out;
SharedReg941_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg941_out;
SharedReg789_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg789_out;
SharedReg400_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg400_out;
SharedReg395_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg395_out;
SharedReg410_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg410_out;
SharedReg395_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg395_out;
SharedReg_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_29_cast <= SharedReg_out;
SharedReg2_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_30_cast <= SharedReg2_out;
SharedReg14_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_31_cast <= SharedReg14_out;
SharedReg4_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_32_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_33_cast <= SharedReg7_out;
SharedReg10_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_34_cast <= SharedReg10_out;
SharedReg9_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_35_cast <= SharedReg9_out;
SharedReg13_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_36_cast <= SharedReg13_out;
SharedReg403_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_37_cast <= SharedReg403_out;
SharedReg400_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_38_cast <= SharedReg400_out;
SharedReg276_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_39_cast <= SharedReg276_out;
SharedReg649_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_40_cast <= SharedReg649_out;
SharedReg4_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_41_cast <= SharedReg4_out;
SharedReg407_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_42_cast <= SharedReg407_out;
SharedReg791_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_43_cast <= SharedReg791_out;
SharedReg797_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_44_cast <= SharedReg797_out;
SharedReg401_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_45_cast <= SharedReg401_out;
SharedReg784_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_46_cast <= SharedReg784_out;
SharedReg395_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_47_cast <= SharedReg395_out;
SharedReg783_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_48_cast <= SharedReg783_out;
SharedReg116_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_49_cast <= SharedReg116_out;
SharedReg531_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_50_cast <= SharedReg531_out;
SharedReg519_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_51_cast <= SharedReg519_out;
SharedReg288_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_52_cast <= SharedReg288_out;
SharedReg395_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_53_cast <= SharedReg395_out;
SharedReg401_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_54_cast <= SharedReg401_out;
SharedReg290_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_55_cast <= SharedReg290_out;
SharedReg783_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_56_cast <= SharedReg783_out;
SharedReg119_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_57_cast <= SharedReg119_out;
SharedReg857_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_58_cast <= SharedReg857_out;
SharedReg663_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_59_cast <= SharedReg663_out;
SharedReg801_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_60_cast <= SharedReg801_out;
SharedReg650_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_61_cast <= SharedReg650_out;
SharedReg649_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_62_cast <= SharedReg649_out;
SharedReg126_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_63_cast <= SharedReg126_out;
SharedReg691_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_64_cast <= SharedReg691_out;
   MUX_Subtract2_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg509_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg398_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg510_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg935_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg265_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg411_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg92_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg118_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg937_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg857_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg397_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg623_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg855_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg267_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg122_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg941_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg789_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg400_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg395_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg410_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg395_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg2_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg696_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg14_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg4_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg7_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg10_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg9_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg13_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg403_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg400_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg276_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg649_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg320_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg4_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg407_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg791_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg797_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg401_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg784_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg395_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg783_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg116_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg531_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg129_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg519_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg288_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg395_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg401_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg290_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg783_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg119_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg857_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg663_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg801_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg932_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg650_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg649_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg126_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg691_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg116_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg128_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg643_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract2_3_impl_0_out);

   Delay1No92_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_3_impl_0_out,
                 Y => Delay1No92_out);

SharedReg514_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg514_out;
SharedReg508_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg508_out;
SharedReg860_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg860_out;
SharedReg855_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg855_out;
SharedReg114_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg114_out;
SharedReg260_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg260_out;
SharedReg658_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg658_out;
SharedReg136_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg136_out;
SharedReg114_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg114_out;
SharedReg953_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg953_out;
SharedReg783_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg783_out;
SharedReg879_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg879_out;
SharedReg137_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg137_out;
SharedReg519_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg519_out;
SharedReg114_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg114_out;
SharedReg114_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg114_out;
SharedReg641_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg641_out;
SharedReg679_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg679_out;
SharedReg503_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg503_out;
SharedReg931_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg931_out;
SharedReg115_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg115_out;
SharedReg114_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg114_out;
SharedReg932_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg932_out;
SharedReg787_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg787_out;
SharedReg516_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg516_out;
SharedReg505_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg505_out;
SharedReg529_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg529_out;
SharedReg787_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg787_out;
SharedReg18_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_29_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_30_cast <= SharedReg20_out;
SharedReg32_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_31_cast <= SharedReg32_out;
SharedReg22_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_32_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_33_cast <= SharedReg25_out;
SharedReg28_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_34_cast <= SharedReg28_out;
SharedReg27_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_35_cast <= SharedReg27_out;
SharedReg31_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_36_cast <= SharedReg31_out;
SharedReg402_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_37_cast <= SharedReg402_out;
SharedReg508_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_38_cast <= SharedReg508_out;
SharedReg127_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_39_cast <= SharedReg127_out;
SharedReg650_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_40_cast <= SharedReg650_out;
SharedReg22_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_41_cast <= SharedReg22_out;
Delay43No10_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_42_cast <= Delay43No10_out;
Delay44No3_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_43_cast <= Delay44No3_out;
SharedReg510_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_44_cast <= SharedReg510_out;
SharedReg503_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_45_cast <= SharedReg503_out;
SharedReg395_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_46_cast <= SharedReg395_out;
SharedReg786_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_47_cast <= SharedReg786_out;
SharedReg403_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_48_cast <= SharedReg403_out;
SharedReg138_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_49_cast <= SharedReg138_out;
SharedReg422_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_50_cast <= SharedReg422_out;
SharedReg803_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_51_cast <= SharedReg803_out;
SharedReg283_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_52_cast <= SharedReg283_out;
SharedReg396_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_53_cast <= SharedReg396_out;
SharedReg395_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_54_cast <= SharedReg395_out;
Delay77No3_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_55_cast <= Delay77No3_out;
SharedReg789_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_56_cast <= SharedReg789_out;
SharedReg261_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_57_cast <= SharedReg261_out;
SharedReg683_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_58_cast <= SharedReg683_out;
SharedReg704_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_59_cast <= SharedReg704_out;
SharedReg811_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_60_cast <= SharedReg811_out;
SharedReg640_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_61_cast <= SharedReg640_out;
SharedReg931_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_62_cast <= SharedReg931_out;
SharedReg115_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_63_cast <= SharedReg115_out;
Delay78No4_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_64_cast <= Delay78No4_out;
   MUX_Subtract2_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg514_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg508_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg783_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg879_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg137_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg519_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg114_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg114_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg641_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg679_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg503_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg931_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg860_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg115_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg114_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg932_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg787_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg516_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg505_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg529_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg787_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg18_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg20_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg855_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg32_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg22_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg25_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg28_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg27_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg31_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg402_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg508_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg127_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg650_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg114_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg22_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => Delay43No10_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => Delay44No3_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg510_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg503_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg395_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg786_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg403_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg138_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg422_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg260_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg803_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg283_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg396_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg395_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => Delay77No3_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg789_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg261_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg683_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg704_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg811_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg658_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg640_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg931_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg115_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => Delay78No4_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg136_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg114_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg953_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract2_3_impl_1_out);

   Delay1No93_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_3_impl_1_out,
                 Y => Delay1No93_out);

Delay1No94_out_to_Subtract2_4_impl_parent_implementedSystem_port_0_cast <= Delay1No94_out;
Delay1No95_out_to_Subtract2_4_impl_parent_implementedSystem_port_1_cast <= Delay1No95_out;
   Subtract2_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_4_impl_out,
                 X => Delay1No94_out_to_Subtract2_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No95_out_to_Subtract2_4_impl_parent_implementedSystem_port_1_cast);

SharedReg801_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg801_out;
SharedReg291_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg291_out;
SharedReg663_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg663_out;
SharedReg687_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg687_out;
SharedReg819_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg819_out;
SharedReg672_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg672_out;
SharedReg865_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg865_out;
SharedReg151_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg151_out;
SharedReg713_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg713_out;
SharedReg525_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg525_out;
SharedReg413_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg413_out;
SharedReg685_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg685_out;
SharedReg717_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg717_out;
SharedReg174_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg174_out;
SharedReg303_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg303_out;
SharedReg856_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg856_out;
SharedReg141_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg141_out;
SharedReg674_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg674_out;
SharedReg664_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg664_out;
SharedReg526_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg526_out;
SharedReg859_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg859_out;
SharedReg290_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg290_out;
SharedReg426_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg426_out;
SharedReg118_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg118_out;
SharedReg142_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg142_out;
SharedReg861_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg861_out;
SharedReg687_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg687_out;
SharedReg412_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg412_out;
SharedReg937_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_29_cast <= SharedReg937_out;
SharedReg292_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_30_cast <= SharedReg292_out;
SharedReg146_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_31_cast <= SharedReg146_out;
SharedReg865_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_32_cast <= SharedReg865_out;
SharedReg807_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_33_cast <= SharedReg807_out;
SharedReg415_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_34_cast <= SharedReg415_out;
SharedReg410_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_35_cast <= SharedReg410_out;
SharedReg425_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_36_cast <= SharedReg425_out;
SharedReg410_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_37_cast <= SharedReg410_out;
SharedReg_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_38_cast <= SharedReg_out;
SharedReg2_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_39_cast <= SharedReg2_out;
SharedReg17_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_40_cast <= SharedReg17_out;
SharedReg695_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_41_cast <= SharedReg695_out;
SharedReg11_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_42_cast <= SharedReg11_out;
SharedReg10_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_43_cast <= SharedReg10_out;
SharedReg9_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_44_cast <= SharedReg9_out;
SharedReg13_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_45_cast <= SharedReg13_out;
SharedReg418_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_46_cast <= SharedReg418_out;
SharedReg415_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_47_cast <= SharedReg415_out;
SharedReg301_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_48_cast <= SharedReg301_out;
SharedReg671_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_49_cast <= SharedReg671_out;
SharedReg4_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_50_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_51_cast <= SharedReg7_out;
SharedReg809_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_52_cast <= SharedReg809_out;
SharedReg815_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_53_cast <= SharedReg815_out;
SharedReg416_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_54_cast <= SharedReg416_out;
SharedReg304_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_55_cast <= SharedReg304_out;
SharedReg873_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_56_cast <= SharedReg873_out;
SharedReg873_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_57_cast <= SharedReg873_out;
SharedReg677_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_58_cast <= SharedReg677_out;
SharedReg831_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_59_cast <= SharedReg831_out;
SharedReg437_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_60_cast <= SharedReg437_out;
SharedReg157_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_61_cast <= SharedReg157_out;
SharedReg665_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_62_cast <= SharedReg665_out;
SharedReg519_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_63_cast <= SharedReg519_out;
SharedReg820_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_64_cast <= SharedReg820_out;
   MUX_Subtract2_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg801_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg291_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg413_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg685_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg717_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg174_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg303_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg856_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg141_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg674_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg664_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg526_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg663_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg859_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg290_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg426_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg118_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg142_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg861_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg687_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg412_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg937_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg292_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg687_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg146_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg865_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg807_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg415_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg410_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg425_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg410_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg2_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg17_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg819_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg695_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg11_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg10_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg9_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg13_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg418_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg415_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg301_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg671_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg4_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg672_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg7_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg809_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg815_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg416_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg304_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg873_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg873_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg677_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg831_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg437_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg865_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg157_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg665_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg519_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg820_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg151_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg713_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg525_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract2_4_impl_0_out);

   Delay1No94_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_4_impl_0_out,
                 Y => Delay1No94_out);

SharedReg807_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg807_out;
SharedReg115_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg115_out;
SharedReg703_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg703_out;
SharedReg727_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg727_out;
SharedReg829_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg829_out;
SharedReg661_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg661_out;
SharedReg855_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg855_out;
SharedReg140_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg140_out;
Delay78No5_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_9_cast <= Delay78No5_out;
SharedReg530_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg530_out;
SharedReg524_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg524_out;
SharedReg690_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg690_out;
SharedReg685_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg685_out;
SharedReg139_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg139_out;
SharedReg285_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg285_out;
SharedReg679_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg679_out;
SharedReg159_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg159_out;
SharedReg855_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg855_out;
SharedReg878_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg878_out;
SharedReg801_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg801_out;
SharedReg702_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg702_out;
SharedReg160_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg160_out;
SharedReg535_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg535_out;
SharedReg139_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg139_out;
SharedReg139_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg139_out;
SharedReg662_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg662_out;
SharedReg723_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg723_out;
SharedReg519_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg519_out;
SharedReg855_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_29_cast <= SharedReg855_out;
SharedReg140_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_30_cast <= SharedReg140_out;
SharedReg139_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_31_cast <= SharedReg139_out;
SharedReg856_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_32_cast <= SharedReg856_out;
SharedReg805_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_33_cast <= SharedReg805_out;
SharedReg532_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_34_cast <= SharedReg532_out;
SharedReg521_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_35_cast <= SharedReg521_out;
SharedReg545_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_36_cast <= SharedReg545_out;
SharedReg805_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_37_cast <= SharedReg805_out;
SharedReg18_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_38_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_39_cast <= SharedReg20_out;
SharedReg35_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_40_cast <= SharedReg35_out;
SharedReg686_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_41_cast <= SharedReg686_out;
SharedReg29_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_42_cast <= SharedReg29_out;
SharedReg28_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_43_cast <= SharedReg28_out;
SharedReg27_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_44_cast <= SharedReg27_out;
SharedReg31_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_45_cast <= SharedReg31_out;
SharedReg417_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_46_cast <= SharedReg417_out;
SharedReg524_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_47_cast <= SharedReg524_out;
SharedReg300_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_48_cast <= SharedReg300_out;
SharedReg672_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_49_cast <= SharedReg672_out;
SharedReg22_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_50_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_51_cast <= SharedReg25_out;
Delay44No4_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_52_cast <= Delay44No4_out;
SharedReg526_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_53_cast <= SharedReg526_out;
SharedReg519_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_54_cast <= SharedReg519_out;
SharedReg114_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_55_cast <= SharedReg114_out;
SharedReg856_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_56_cast <= SharedReg856_out;
SharedReg642_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_57_cast <= SharedReg642_out;
SharedReg720_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_58_cast <= SharedReg720_out;
SharedReg834_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_59_cast <= SharedReg834_out;
Delay43No12_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_60_cast <= Delay43No12_out;
SharedReg291_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_61_cast <= SharedReg291_out;
Delay76No4_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_62_cast <= Delay76No4_out;
SharedReg806_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_63_cast <= SharedReg806_out;
SharedReg425_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_64_cast <= SharedReg425_out;
   MUX_Subtract2_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg807_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg115_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg524_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg690_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg685_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg139_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg285_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg679_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg159_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg855_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg878_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg801_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg703_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg702_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg160_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg535_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg139_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg139_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg662_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg723_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg519_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg855_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg140_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg727_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg139_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg856_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg805_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg532_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg521_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg545_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg805_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg18_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg20_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg35_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg829_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg686_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg29_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg28_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg27_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg31_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg417_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg524_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg300_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg672_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg22_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg661_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg25_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => Delay44No4_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg526_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg519_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg114_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg856_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg642_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg720_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg834_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => Delay43No12_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg855_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg291_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => Delay76No4_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg806_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg425_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg140_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay78No5_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg530_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract2_4_impl_1_out);

   Delay1No95_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_4_impl_1_out,
                 Y => Delay1No95_out);

Delay1No96_out_to_Subtract2_5_impl_parent_implementedSystem_port_0_cast <= Delay1No96_out;
Delay1No97_out_to_Subtract2_5_impl_parent_implementedSystem_port_1_cast <= Delay1No97_out;
   Subtract2_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_5_impl_out,
                 X => Delay1No96_out_to_Subtract2_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No97_out_to_Subtract2_5_impl_parent_implementedSystem_port_1_cast);

SharedReg425_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg425_out;
SharedReg819_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg819_out;
SharedReg141_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg141_out;
SharedReg997_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg997_out;
SharedReg563_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg563_out;
SharedReg166_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg166_out;
SharedReg425_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg425_out;
SharedReg431_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg431_out;
SharedReg168_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg168_out;
SharedReg538_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg538_out;
SharedReg535_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg535_out;
SharedReg163_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg163_out;
SharedReg985_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg985_out;
SharedReg188_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_14_cast <= SharedReg188_out;
SharedReg163_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_15_cast <= SharedReg163_out;
SharedReg320_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_16_cast <= SharedReg320_out;
SharedReg687_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_17_cast <= SharedReg687_out;
SharedReg446_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_18_cast <= SharedReg446_out;
SharedReg429_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_19_cast <= SharedReg429_out;
SharedReg539_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_20_cast <= SharedReg539_out;
SharedReg538_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_21_cast <= SharedReg538_out;
SharedReg882_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_22_cast <= SharedReg882_out;
SharedReg440_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_23_cast <= SharedReg440_out;
SharedReg820_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_24_cast <= SharedReg820_out;
SharedReg871_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_25_cast <= SharedReg871_out;
SharedReg426_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_26_cast <= SharedReg426_out;
SharedReg884_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_27_cast <= SharedReg884_out;
SharedReg313_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_28_cast <= SharedReg313_out;
SharedReg425_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_29_cast <= SharedReg425_out;
SharedReg168_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_30_cast <= SharedReg168_out;
SharedReg425_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_31_cast <= SharedReg425_out;
SharedReg427_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_32_cast <= SharedReg427_out;
SharedReg535_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_33_cast <= SharedReg535_out;
SharedReg667_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_34_cast <= SharedReg667_out;
SharedReg427_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_35_cast <= SharedReg427_out;
SharedReg441_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_36_cast <= SharedReg441_out;
SharedReg801_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_37_cast <= SharedReg801_out;
SharedReg1_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1_out;
SharedReg3_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_39_cast <= SharedReg3_out;
SharedReg172_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_40_cast <= SharedReg172_out;
SharedReg440_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_41_cast <= SharedReg440_out;
SharedReg825_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_42_cast <= SharedReg825_out;
SharedReg12_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_43_cast <= SharedReg12_out;
SharedReg16_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_44_cast <= SharedReg16_out;
SharedReg425_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_45_cast <= SharedReg425_out;
SharedReg525_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_46_cast <= SharedReg525_out;
SharedReg522_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_47_cast <= SharedReg522_out;
SharedReg146_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_48_cast <= SharedReg146_out;
SharedReg14_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_49_cast <= SharedReg14_out;
SharedReg6_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_50_cast <= SharedReg6_out;
SharedReg11_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_51_cast <= SharedReg11_out;
SharedReg522_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_52_cast <= SharedReg522_out;
SharedReg419_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_53_cast <= SharedReg419_out;
SharedReg8_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_54_cast <= SharedReg8_out;
SharedReg433_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_55_cast <= SharedReg433_out;
SharedReg430_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_56_cast <= SharedReg430_out;
SharedReg324_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_57_cast <= SharedReg324_out;
SharedReg716_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_58_cast <= SharedReg716_out;
SharedReg14_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_59_cast <= SharedReg14_out;
SharedReg4_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_60_cast <= SharedReg4_out;
SharedReg827_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_61_cast <= SharedReg827_out;
SharedReg833_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_62_cast <= SharedReg833_out;
SharedReg431_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_63_cast <= SharedReg431_out;
SharedReg326_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_64_cast <= SharedReg326_out;
   MUX_Subtract2_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg425_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg819_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg535_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg163_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg985_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg188_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg163_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg320_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg687_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg446_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg429_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg539_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg141_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg538_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg882_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg440_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg820_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg871_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg426_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg884_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg313_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg425_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg168_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg997_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg425_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg427_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg535_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg667_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg427_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg441_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg801_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg3_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg172_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg563_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg440_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg825_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg12_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg16_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg425_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg525_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg522_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg146_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg14_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg6_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg166_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg11_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg522_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg419_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg8_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg433_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg430_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg324_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg716_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg14_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg4_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg425_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg827_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg833_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg431_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg326_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg431_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg168_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg538_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract2_5_impl_0_out);

   Delay1No96_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_5_impl_0_out,
                 Y => Delay1No96_out);

SharedReg822_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg822_out;
SharedReg433_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg433_out;
SharedReg330_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg330_out;
SharedReg996_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg996_out;
SharedReg452_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg452_out;
SharedReg162_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg162_out;
SharedReg426_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg426_out;
SharedReg425_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg425_out;
Delay77No5_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_9_cast <= Delay77No5_out;
SharedReg535_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg535_out;
SharedReg821_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg821_out;
SharedReg169_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg169_out;
SharedReg904_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg904_out;
SharedReg206_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_14_cast <= SharedReg206_out;
SharedReg165_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_15_cast <= SharedReg165_out;
SharedReg310_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_16_cast <= SharedReg310_out;
SharedReg711_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_17_cast <= SharedReg711_out;
SharedReg440_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_18_cast <= SharedReg440_out;
SharedReg835_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_19_cast <= SharedReg835_out;
SharedReg826_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_20_cast <= SharedReg826_out;
SharedReg824_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_21_cast <= SharedReg824_out;
SharedReg712_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_22_cast <= SharedReg712_out;
SharedReg450_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_23_cast <= SharedReg450_out;
SharedReg535_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_24_cast <= SharedReg535_out;
SharedReg708_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_25_cast <= SharedReg708_out;
SharedReg535_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_26_cast <= SharedReg535_out;
SharedReg711_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_27_cast <= SharedReg711_out;
SharedReg329_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_28_cast <= SharedReg329_out;
SharedReg536_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_29_cast <= SharedReg536_out;
SharedReg183_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_30_cast <= SharedReg183_out;
SharedReg820_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_31_cast <= SharedReg820_out;
SharedReg535_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_32_cast <= SharedReg535_out;
SharedReg828_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_33_cast <= SharedReg828_out;
SharedReg685_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_34_cast <= SharedReg685_out;
SharedReg822_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_35_cast <= SharedReg822_out;
SharedReg551_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_36_cast <= SharedReg551_out;
SharedReg804_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_37_cast <= SharedReg804_out;
SharedReg19_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_38_cast <= SharedReg19_out;
SharedReg21_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_39_cast <= SharedReg21_out;
SharedReg163_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_40_cast <= SharedReg163_out;
SharedReg838_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_41_cast <= SharedReg838_out;
SharedReg823_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_42_cast <= SharedReg823_out;
SharedReg30_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_43_cast <= SharedReg30_out;
SharedReg34_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_44_cast <= SharedReg34_out;
SharedReg537_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_45_cast <= SharedReg537_out;
SharedReg807_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_46_cast <= SharedReg807_out;
SharedReg807_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_47_cast <= SharedReg807_out;
SharedReg147_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_48_cast <= SharedReg147_out;
SharedReg32_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_49_cast <= SharedReg32_out;
SharedReg24_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_50_cast <= SharedReg24_out;
SharedReg29_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_51_cast <= SharedReg29_out;
SharedReg801_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_52_cast <= SharedReg801_out;
SharedReg417_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_53_cast <= SharedReg417_out;
SharedReg26_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_54_cast <= SharedReg26_out;
SharedReg432_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_55_cast <= SharedReg432_out;
SharedReg540_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_56_cast <= SharedReg540_out;
SharedReg323_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_57_cast <= SharedReg323_out;
SharedReg696_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_58_cast <= SharedReg696_out;
SharedReg32_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_59_cast <= SharedReg32_out;
SharedReg22_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_60_cast <= SharedReg22_out;
Delay44No5_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_61_cast <= Delay44No5_out;
SharedReg542_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_62_cast <= SharedReg542_out;
SharedReg535_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_63_cast <= SharedReg535_out;
SharedReg285_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_64_cast <= SharedReg285_out;
   MUX_Subtract2_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg822_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg433_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg821_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg169_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg904_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg206_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg165_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg310_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg711_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg440_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg835_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg826_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg330_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg824_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg712_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg450_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg535_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg708_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg535_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg711_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg329_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg536_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg183_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg996_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg820_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg535_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg828_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg685_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg822_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg551_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg804_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg19_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg21_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg163_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg452_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg838_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg823_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg30_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg34_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg537_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg807_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg807_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg147_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg32_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg24_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg162_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg29_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg801_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg417_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg26_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg432_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg540_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg323_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg696_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg32_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg22_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg426_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => Delay44No5_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg542_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg535_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg285_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg425_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay77No5_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg535_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract2_5_impl_1_out);

   Delay1No97_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_5_impl_1_out,
                 Y => Delay1No97_out);

Delay1No98_out_to_Subtract2_6_impl_parent_implementedSystem_port_0_cast <= Delay1No98_out;
Delay1No99_out_to_Subtract2_6_impl_parent_implementedSystem_port_1_cast <= Delay1No99_out;
   Subtract2_6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_6_impl_out,
                 X => Delay1No98_out_to_Subtract2_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No99_out_to_Subtract2_6_impl_parent_implementedSystem_port_1_cast);

SharedReg6_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg6_out;
SharedReg_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg_out;
SharedReg2_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg2_out;
SharedReg2_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg2_out;
SharedReg8_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg8_out;
SharedReg9_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg9_out;
SharedReg9_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg9_out;
SharedReg10_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg10_out;
SharedReg13_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg13_out;
SharedReg17_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg17_out;
SharedReg17_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg17_out;
SharedReg699_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg699_out;
SharedReg446_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_13_cast <= SharedReg446_out;
SharedReg696_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_14_cast <= SharedReg696_out;
SharedReg322_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_15_cast <= SharedReg322_out;
SharedReg200_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_16_cast <= SharedReg200_out;
SharedReg695_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_17_cast <= SharedReg695_out;
SharedReg325_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_18_cast <= SharedReg325_out;
SharedReg332_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_19_cast <= SharedReg332_out;
SharedReg837_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_20_cast <= SharedReg837_out;
SharedReg442_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_21_cast <= SharedReg442_out;
SharedReg195_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_22_cast <= SharedReg195_out;
SharedReg142_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_23_cast <= SharedReg142_out;
SharedReg695_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_24_cast <= SharedReg695_out;
SharedReg201_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_25_cast <= SharedReg201_out;
SharedReg427_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_26_cast <= SharedReg427_out;
SharedReg172_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_27_cast <= SharedReg172_out;
SharedReg430_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_28_cast <= SharedReg430_out;
SharedReg993_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_29_cast <= SharedReg993_out;
SharedReg168_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_30_cast <= SharedReg168_out;
SharedReg691_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_31_cast <= SharedReg691_out;
SharedReg442_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_32_cast <= SharedReg442_out;
SharedReg180_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_33_cast <= SharedReg180_out;
SharedReg699_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_34_cast <= SharedReg699_out;
SharedReg316_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_35_cast <= SharedReg316_out;
SharedReg861_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_36_cast <= SharedReg861_out;
SharedReg849_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_37_cast <= SharedReg849_out;
SharedReg542_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_38_cast <= SharedReg542_out;
SharedReg334_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_39_cast <= SharedReg334_out;
SharedReg689_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_40_cast <= SharedReg689_out;
SharedReg434_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_41_cast <= SharedReg434_out;
SharedReg541_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_42_cast <= SharedReg541_out;
SharedReg165_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_43_cast <= SharedReg165_out;
SharedReg334_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_44_cast <= SharedReg334_out;
SharedReg686_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_45_cast <= SharedReg686_out;
SharedReg538_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_46_cast <= SharedReg538_out;
SharedReg425_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_47_cast <= SharedReg425_out;
SharedReg819_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_48_cast <= SharedReg819_out;
SharedReg884_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_49_cast <= SharedReg884_out;
SharedReg425_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_50_cast <= SharedReg425_out;
SharedReg337_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_51_cast <= SharedReg337_out;
SharedReg428_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_52_cast <= SharedReg428_out;
SharedReg710_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_53_cast <= SharedReg710_out;
SharedReg315_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_54_cast <= SharedReg315_out;
SharedReg191_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_55_cast <= SharedReg191_out;
SharedReg689_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_56_cast <= SharedReg689_out;
SharedReg551_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_57_cast <= SharedReg551_out;
SharedReg541_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_58_cast <= SharedReg541_out;
SharedReg538_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_59_cast <= SharedReg538_out;
SharedReg535_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_60_cast <= SharedReg535_out;
SharedReg551_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_61_cast <= SharedReg551_out;
SharedReg143_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_62_cast <= SharedReg143_out;
SharedReg994_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_63_cast <= SharedReg994_out;
   MUX_Subtract2_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_63_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg6_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg17_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg699_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg446_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg696_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg322_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg200_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg695_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg325_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg332_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg837_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg2_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg442_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg195_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg142_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg695_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg201_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg427_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg172_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg430_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg993_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg168_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg2_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg691_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg442_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg180_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg699_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg316_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg861_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg849_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg542_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg334_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg689_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg8_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg434_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg541_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg165_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg334_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg686_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg538_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg425_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg819_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg884_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg425_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg9_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg337_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg428_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg710_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg315_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg191_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg689_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg551_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg541_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg538_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg535_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg9_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg551_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg143_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg994_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_63_cast,
                 iS_7 => SharedReg10_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg13_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg17_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Subtract2_6_impl_0_LUT_out,
                 oMux => MUX_Subtract2_6_impl_0_out);

   Delay1No98_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_6_impl_0_out,
                 Y => Delay1No98_out);

SharedReg18_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg20_out;
SharedReg20_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg20_out;
SharedReg24_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg24_out;
SharedReg26_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg26_out;
SharedReg27_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg27_out;
SharedReg27_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg27_out;
SharedReg28_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg28_out;
SharedReg31_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg31_out;
SharedReg35_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg35_out;
SharedReg35_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg35_out;
SharedReg551_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg551_out;
SharedReg140_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_13_cast <= SharedReg140_out;
SharedReg685_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_14_cast <= SharedReg685_out;
SharedReg310_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_15_cast <= SharedReg310_out;
SharedReg338_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_16_cast <= SharedReg338_out;
SharedReg448_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_17_cast <= SharedReg448_out;
SharedReg551_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_18_cast <= SharedReg551_out;
SharedReg343_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_19_cast <= SharedReg343_out;
SharedReg535_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_20_cast <= SharedReg535_out;
SharedReg310_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_21_cast <= SharedReg310_out;
SharedReg548_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_22_cast <= SharedReg548_out;
SharedReg857_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_23_cast <= SharedReg857_out;
SharedReg852_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_24_cast <= SharedReg852_out;
SharedReg662_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_25_cast <= SharedReg662_out;
SharedReg332_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_26_cast <= SharedReg332_out;
SharedReg840_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_27_cast <= SharedReg840_out;
SharedReg708_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_28_cast <= SharedReg708_out;
SharedReg143_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_29_cast <= SharedReg143_out;
SharedReg164_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_30_cast <= SharedReg164_out;
SharedReg685_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_31_cast <= SharedReg685_out;
SharedReg819_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_32_cast <= SharedReg819_out;
SharedReg318_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_33_cast <= SharedReg318_out;
SharedReg994_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_34_cast <= SharedReg994_out;
SharedReg163_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_35_cast <= SharedReg163_out;
SharedReg708_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_36_cast <= SharedReg708_out;
SharedReg206_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_37_cast <= SharedReg206_out;
SharedReg432_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_38_cast <= SharedReg432_out;
SharedReg706_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_39_cast <= SharedReg706_out;
SharedReg825_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_40_cast <= SharedReg825_out;
SharedReg182_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_41_cast <= SharedReg182_out;
SharedReg347_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_42_cast <= SharedReg347_out;
SharedReg825_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_43_cast <= SharedReg825_out;
SharedReg1001_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_44_cast <= SharedReg1001_out;
SharedReg537_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_45_cast <= SharedReg537_out;
SharedReg723_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_46_cast <= SharedReg723_out;
SharedReg825_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_47_cast <= SharedReg825_out;
SharedReg707_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_48_cast <= SharedReg707_out;
SharedReg823_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_49_cast <= SharedReg823_out;
SharedReg540_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_50_cast <= SharedReg540_out;
SharedReg183_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_51_cast <= SharedReg183_out;
SharedReg903_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_52_cast <= SharedReg903_out;
SharedReg701_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_53_cast <= SharedReg701_out;
SharedReg183_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_54_cast <= SharedReg183_out;
SharedReg348_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_55_cast <= SharedReg348_out;
SharedReg164_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_56_cast <= SharedReg164_out;
SharedReg187_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_57_cast <= SharedReg187_out;
SharedReg839_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_58_cast <= SharedReg839_out;
SharedReg685_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_59_cast <= SharedReg685_out;
SharedReg546_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_60_cast <= SharedReg546_out;
SharedReg824_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_61_cast <= SharedReg824_out;
SharedReg842_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_62_cast <= SharedReg842_out;
SharedReg819_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_63_cast <= SharedReg819_out;
   MUX_Subtract2_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_63_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg18_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg20_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg35_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg551_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg140_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg685_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg310_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg338_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg448_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg551_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg343_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg535_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg20_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg310_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg548_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg857_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg852_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg662_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg332_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg840_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg708_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg143_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg164_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg24_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg685_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg819_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg318_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg994_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg163_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg708_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg206_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg432_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg706_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg825_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg26_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg182_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg347_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg825_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1001_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg537_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg723_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg825_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg707_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg823_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg540_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg27_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg183_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg903_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg701_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg183_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg348_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg164_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg187_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg839_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg685_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg546_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg27_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg824_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg842_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg819_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_63_cast,
                 iS_7 => SharedReg28_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg31_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg35_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Subtract2_6_impl_1_LUT_out,
                 oMux => MUX_Subtract2_6_impl_1_out);

   Delay1No99_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_6_impl_1_out,
                 Y => Delay1No99_out);

Delay1No100_out_to_Product32_0_impl_parent_implementedSystem_port_0_cast <= Delay1No100_out;
Delay1No101_out_to_Product32_0_impl_parent_implementedSystem_port_1_cast <= Delay1No101_out;
   Product32_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_0_impl_out,
                 X => Delay1No100_out_to_Product32_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No101_out_to_Product32_0_impl_parent_implementedSystem_port_1_cast);

SharedReg568_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg568_out;
SharedReg1134_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1134_out;
SharedReg1149_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1149_out;
SharedReg1055_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1055_out;
SharedReg1056_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1056_out;
SharedReg36_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg36_out;
SharedReg957_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg957_out;
SharedReg1170_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1170_out;
SharedReg36_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg36_out;
SharedReg1005_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1005_out;
SharedReg1059_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1059_out;
SharedReg961_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg961_out;
SharedReg213_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg213_out;
SharedReg1109_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1109_out;
SharedReg1009_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1009_out;
SharedReg1169_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1169_out;
SharedReg1167_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1167_out;
SharedReg217_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg217_out;
SharedReg43_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg43_out;
SharedReg1012_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1012_out;
SharedReg1065_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1065_out;
SharedReg1122_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1122_out;
SharedReg1014_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1014_out;
SharedReg220_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg220_out;
SharedReg1016_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1016_out;
SharedReg1068_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1068_out;
SharedReg1069_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1069_out;
SharedReg577_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg577_out;
SharedReg1097_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1097_out;
SharedReg1098_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1098_out;
SharedReg971_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_31_cast <= SharedReg971_out;
SharedReg1100_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1100_out;
SharedReg966_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_33_cast <= SharedReg966_out;
SharedReg1053_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1053_out;
SharedReg1102_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1102_out;
SharedReg1162_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1162_out;
SharedReg1116_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1116_out;
SharedReg1110_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1110_out;
SharedReg567_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_39_cast <= SharedReg567_out;
SharedReg1118_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1118_out;
SharedReg1112_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1112_out;
SharedReg1157_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1157_out;
SharedReg1026_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1026_out;
SharedReg965_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_44_cast <= SharedReg965_out;
SharedReg572_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_45_cast <= SharedReg572_out;
SharedReg1078_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1078_out;
SharedReg44_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_47_cast <= SharedReg44_out;
SharedReg1165_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1165_out;
SharedReg574_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_49_cast <= SharedReg574_out;
SharedReg1139_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1139_out;
SharedReg1126_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1126_out;
SharedReg1127_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1127_out;
SharedReg962_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_53_cast <= SharedReg962_out;
SharedReg1141_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1141_out;
SharedReg1128_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1128_out;
SharedReg1054_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1054_out;
SharedReg957_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_57_cast <= SharedReg957_out;
SharedReg957_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_58_cast <= SharedReg957_out;
SharedReg1129_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1129_out;
SharedReg1144_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1144_out;
SharedReg1130_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1130_out;
SharedReg1131_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1131_out;
SharedReg1146_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1146_out;
SharedReg568_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_64_cast <= SharedReg568_out;
   MUX_Product32_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg568_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1134_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1059_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg961_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg213_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1109_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1009_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1169_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1167_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg217_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg43_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1012_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1149_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1065_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1122_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1014_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg220_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1016_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1068_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1069_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg577_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1097_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1098_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1055_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg971_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1100_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg966_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1053_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1102_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1162_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1116_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1110_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg567_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1118_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1056_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1112_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1157_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1026_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg965_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg572_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1078_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg44_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1165_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg574_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1139_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg36_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1126_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1127_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg962_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1141_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1128_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1054_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg957_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg957_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1129_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1144_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg957_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1130_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1131_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1146_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg568_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1170_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg36_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1005_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product32_0_impl_0_out);

   Delay1No100_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_0_impl_0_out,
                 Y => Delay1No100_out);

SharedReg1148_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1148_out;
SharedReg569_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg569_out;
SharedReg569_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg569_out;
SharedReg979_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg979_out;
SharedReg976_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg976_out;
SharedReg1095_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1095_out;
SharedReg1057_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1057_out;
SharedReg957_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg957_out;
SharedReg1058_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1058_out;
SharedReg208_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg208_out;
SharedReg37_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg37_out;
SharedReg1171_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1171_out;
SharedReg1060_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1060_out;
SharedReg571_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg571_out;
SharedReg965_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg965_out;
SharedReg960_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg960_out;
SharedReg961_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg961_out;
SharedReg1063_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1063_out;
SharedReg1064_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1064_out;
SharedReg579_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg579_out;
SharedReg46_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg46_out;
SharedReg577_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg577_out;
SharedReg222_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg222_out;
SharedReg1066_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1066_out;
SharedReg48_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg48_out;
SharedReg223_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg223_out;
SharedReg49_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg49_out;
SharedReg1096_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1096_out;
SharedReg47_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_29_cast <= SharedReg47_out;
SharedReg578_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_30_cast <= SharedReg578_out;
SharedReg1099_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_31_cast <= SharedReg1099_out;
SharedReg971_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_32_cast <= SharedReg971_out;
SharedReg1101_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_33_cast <= SharedReg1101_out;
SharedReg967_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_34_cast <= SharedReg967_out;
SharedReg217_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_35_cast <= SharedReg217_out;
SharedReg567_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_36_cast <= SharedReg567_out;
SharedReg957_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_37_cast <= SharedReg957_out;
SharedReg958_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_38_cast <= SharedReg958_out;
SharedReg1163_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_39_cast <= SharedReg1163_out;
SharedReg957_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_40_cast <= SharedReg957_out;
SharedReg958_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_41_cast <= SharedReg958_out;
SharedReg570_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_42_cast <= SharedReg570_out;
SharedReg40_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_43_cast <= SharedReg40_out;
SharedReg1164_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_44_cast <= SharedReg1164_out;
SharedReg1077_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_45_cast <= SharedReg1077_out;
SharedReg964_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_46_cast <= SharedReg964_out;
SharedReg1079_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_47_cast <= SharedReg1079_out;
SharedReg574_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_48_cast <= SharedReg574_out;
SharedReg1138_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_49_cast <= SharedReg1138_out;
SharedReg965_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_50_cast <= SharedReg965_out;
SharedReg966_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_51_cast <= SharedReg966_out;
SharedReg961_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_52_cast <= SharedReg961_out;
SharedReg1140_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_53_cast <= SharedReg1140_out;
SharedReg572_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_54_cast <= SharedReg572_out;
SharedReg573_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_55_cast <= SharedReg573_out;
SharedReg226_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_56_cast <= SharedReg226_out;
SharedReg1142_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1142_out;
SharedReg1143_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_58_cast <= SharedReg1143_out;
SharedReg958_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_59_cast <= SharedReg958_out;
SharedReg958_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_60_cast <= SharedReg958_out;
SharedReg959_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_61_cast <= SharedReg959_out;
SharedReg962_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_62_cast <= SharedReg962_out;
SharedReg568_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_63_cast <= SharedReg568_out;
SharedReg1147_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_64_cast <= SharedReg1147_out;
   MUX_Product32_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1148_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg569_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg37_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1171_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1060_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg571_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg965_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg960_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg961_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1063_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1064_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg579_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg569_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg46_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg577_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg222_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1066_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg48_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg223_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg49_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1096_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg47_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg578_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg979_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1099_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg971_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1101_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg967_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg217_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg567_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg957_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg958_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1163_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg957_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg976_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg958_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg570_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg40_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1164_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1077_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg964_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1079_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg574_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1138_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg965_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1095_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg966_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg961_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1140_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg572_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg573_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg226_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1142_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1143_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg958_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg958_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1057_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg959_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg962_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg568_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1147_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg957_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1058_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg208_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product32_0_impl_1_out);

   Delay1No101_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_0_impl_1_out,
                 Y => Delay1No101_out);

Delay1No102_out_to_Product32_1_impl_parent_implementedSystem_port_0_cast <= Delay1No102_out;
Delay1No103_out_to_Product32_1_impl_parent_implementedSystem_port_1_cast <= Delay1No103_out;
   Product32_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_1_impl_out,
                 X => Delay1No102_out_to_Product32_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No103_out_to_Product32_1_impl_parent_implementedSystem_port_1_cast);

SharedReg1054_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1054_out;
SharedReg593_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg593_out;
SharedReg593_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg593_out;
SharedReg1129_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1129_out;
SharedReg1144_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1144_out;
SharedReg1130_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1130_out;
SharedReg1131_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1131_out;
SharedReg1146_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1146_out;
SharedReg594_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg594_out;
SharedReg594_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg594_out;
SharedReg1134_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1134_out;
SharedReg1149_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1149_out;
SharedReg1055_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1055_out;
SharedReg1056_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1056_out;
SharedReg62_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg62_out;
SharedReg906_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg906_out;
SharedReg1170_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1170_out;
SharedReg62_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg62_out;
SharedReg1005_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1005_out;
SharedReg1059_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1059_out;
SharedReg910_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg910_out;
SharedReg239_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg239_out;
SharedReg1109_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1109_out;
SharedReg1009_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1009_out;
SharedReg1169_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1169_out;
SharedReg1167_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1167_out;
SharedReg243_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg243_out;
SharedReg69_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg69_out;
SharedReg1012_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1012_out;
SharedReg1065_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1065_out;
SharedReg1122_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1122_out;
SharedReg1014_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1014_out;
SharedReg246_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_33_cast <= SharedReg246_out;
SharedReg1016_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1016_out;
SharedReg1068_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1068_out;
SharedReg1069_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1069_out;
SharedReg603_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_37_cast <= SharedReg603_out;
SharedReg1097_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1097_out;
SharedReg1098_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1098_out;
SharedReg919_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_40_cast <= SharedReg919_out;
SharedReg1100_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1100_out;
SharedReg915_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_42_cast <= SharedReg915_out;
SharedReg1053_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1053_out;
SharedReg1102_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1102_out;
SharedReg1162_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1162_out;
SharedReg1116_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1116_out;
SharedReg1110_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1110_out;
SharedReg593_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_48_cast <= SharedReg593_out;
SharedReg1118_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1118_out;
SharedReg1112_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1112_out;
SharedReg1157_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1157_out;
SharedReg1026_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1026_out;
SharedReg601_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_53_cast <= SharedReg601_out;
SharedReg598_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_54_cast <= SharedReg598_out;
SharedReg1078_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1078_out;
SharedReg70_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_56_cast <= SharedReg70_out;
SharedReg1165_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1165_out;
SharedReg600_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_58_cast <= SharedReg600_out;
SharedReg1139_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1139_out;
SharedReg1126_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1126_out;
SharedReg1127_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1127_out;
SharedReg911_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_62_cast <= SharedReg911_out;
SharedReg1141_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1141_out;
SharedReg1128_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1128_out;
   MUX_Product32_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1054_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg593_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1134_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1149_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1055_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1056_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg62_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg906_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1170_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg62_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1005_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1059_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg593_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg910_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg239_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1109_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1009_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1169_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1167_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg243_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg69_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1012_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1065_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1129_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1122_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1014_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg246_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1016_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1068_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1069_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg603_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1097_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1098_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg919_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1144_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1100_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg915_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1053_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1102_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1162_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1116_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1110_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg593_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1118_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1112_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1130_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1157_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1026_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg601_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg598_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1078_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg70_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1165_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg600_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1139_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1126_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1131_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1127_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg911_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1141_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1128_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1146_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg594_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg594_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product32_1_impl_0_out);

   Delay1No102_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_1_impl_0_out,
                 Y => Delay1No102_out);

SharedReg252_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg252_out;
SharedReg1142_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1142_out;
SharedReg1143_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1143_out;
SharedReg594_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg594_out;
SharedReg594_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg594_out;
SharedReg595_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg595_out;
SharedReg598_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg598_out;
SharedReg594_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg594_out;
SharedReg1147_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1147_out;
SharedReg1148_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1148_out;
SharedReg595_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg595_out;
SharedReg595_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg595_out;
SharedReg927_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg927_out;
SharedReg924_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg924_out;
SharedReg1095_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1095_out;
SharedReg1057_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1057_out;
SharedReg906_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg906_out;
SharedReg1058_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1058_out;
SharedReg234_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg234_out;
SharedReg63_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg63_out;
SharedReg1171_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1171_out;
SharedReg1060_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1060_out;
SharedReg597_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg597_out;
SharedReg914_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg914_out;
SharedReg909_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg909_out;
SharedReg910_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg910_out;
SharedReg1063_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1063_out;
SharedReg1064_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1064_out;
SharedReg605_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_29_cast <= SharedReg605_out;
SharedReg72_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_30_cast <= SharedReg72_out;
SharedReg603_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_31_cast <= SharedReg603_out;
SharedReg248_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_32_cast <= SharedReg248_out;
SharedReg1066_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_33_cast <= SharedReg1066_out;
SharedReg74_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_34_cast <= SharedReg74_out;
SharedReg249_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_35_cast <= SharedReg249_out;
SharedReg75_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_36_cast <= SharedReg75_out;
SharedReg1096_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_37_cast <= SharedReg1096_out;
SharedReg73_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_38_cast <= SharedReg73_out;
SharedReg604_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_39_cast <= SharedReg604_out;
SharedReg1099_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_40_cast <= SharedReg1099_out;
SharedReg919_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_41_cast <= SharedReg919_out;
SharedReg1101_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_42_cast <= SharedReg1101_out;
SharedReg916_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_43_cast <= SharedReg916_out;
SharedReg243_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_44_cast <= SharedReg243_out;
SharedReg957_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_45_cast <= SharedReg957_out;
SharedReg957_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_46_cast <= SharedReg957_out;
SharedReg958_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_47_cast <= SharedReg958_out;
SharedReg1163_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_48_cast <= SharedReg1163_out;
SharedReg906_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_49_cast <= SharedReg906_out;
SharedReg907_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_50_cast <= SharedReg907_out;
SharedReg596_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_51_cast <= SharedReg596_out;
SharedReg66_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_52_cast <= SharedReg66_out;
SharedReg1164_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_53_cast <= SharedReg1164_out;
SharedReg1077_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_54_cast <= SharedReg1077_out;
SharedReg913_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_55_cast <= SharedReg913_out;
SharedReg1079_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_56_cast <= SharedReg1079_out;
SharedReg600_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_57_cast <= SharedReg600_out;
SharedReg1138_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_58_cast <= SharedReg1138_out;
SharedReg914_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_59_cast <= SharedReg914_out;
SharedReg915_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_60_cast <= SharedReg915_out;
SharedReg910_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_61_cast <= SharedReg910_out;
SharedReg1140_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_62_cast <= SharedReg1140_out;
SharedReg598_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_63_cast <= SharedReg598_out;
SharedReg599_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_64_cast <= SharedReg599_out;
   MUX_Product32_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg252_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1142_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg595_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg595_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg927_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg924_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1095_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1057_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg906_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1058_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg234_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg63_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1143_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1171_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1060_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg597_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg914_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg909_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg910_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1063_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1064_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg605_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg72_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg594_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg603_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg248_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1066_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg74_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg249_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg75_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1096_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg73_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg604_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1099_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg594_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg919_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1101_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg916_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg243_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg957_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg957_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg958_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1163_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg906_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg907_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg595_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg596_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg66_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1164_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1077_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg913_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1079_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg600_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1138_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg914_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg915_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg598_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg910_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1140_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg598_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg599_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg594_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1147_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1148_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product32_1_impl_1_out);

   Delay1No103_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_1_impl_1_out,
                 Y => Delay1No103_out);

Delay1No104_out_to_Product32_2_impl_parent_implementedSystem_port_0_cast <= Delay1No104_out;
Delay1No105_out_to_Product32_2_impl_parent_implementedSystem_port_1_cast <= Delay1No105_out;
   Product32_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_2_impl_out,
                 X => Delay1No104_out_to_Product32_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No105_out_to_Product32_2_impl_parent_implementedSystem_port_1_cast);

SharedReg95_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg95_out;
SharedReg1165_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1165_out;
SharedReg913_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg913_out;
SharedReg1139_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1139_out;
SharedReg1126_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1126_out;
SharedReg1127_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1127_out;
SharedReg622_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg622_out;
SharedReg1141_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1141_out;
SharedReg1128_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1128_out;
SharedReg1054_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1054_out;
SharedReg617_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg617_out;
SharedReg617_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg617_out;
SharedReg1129_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1129_out;
SharedReg1144_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1144_out;
SharedReg1130_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1130_out;
SharedReg1131_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1131_out;
SharedReg1146_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1146_out;
SharedReg618_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg618_out;
SharedReg618_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg618_out;
SharedReg1134_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1134_out;
SharedReg1149_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1149_out;
SharedReg1055_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1055_out;
SharedReg1056_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1056_out;
SharedReg88_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg88_out;
SharedReg931_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg931_out;
SharedReg1170_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1170_out;
SharedReg88_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg88_out;
SharedReg1005_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1005_out;
SharedReg1059_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1059_out;
SharedReg935_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_30_cast <= SharedReg935_out;
SharedReg265_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_31_cast <= SharedReg265_out;
SharedReg1109_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1109_out;
SharedReg1009_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1009_out;
SharedReg1169_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1169_out;
SharedReg1167_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1167_out;
SharedReg269_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_36_cast <= SharedReg269_out;
SharedReg94_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_37_cast <= SharedReg94_out;
SharedReg1012_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1012_out;
SharedReg1065_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1065_out;
SharedReg1122_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1122_out;
SharedReg1014_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1014_out;
SharedReg272_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_42_cast <= SharedReg272_out;
SharedReg1016_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1016_out;
SharedReg1068_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1068_out;
SharedReg1069_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1069_out;
SharedReg628_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_46_cast <= SharedReg628_out;
SharedReg1097_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1097_out;
SharedReg1098_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1098_out;
SharedReg944_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_49_cast <= SharedReg944_out;
SharedReg1100_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1100_out;
SharedReg940_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_51_cast <= SharedReg940_out;
SharedReg1053_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1053_out;
SharedReg1102_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1102_out;
SharedReg1162_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1162_out;
SharedReg1116_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1116_out;
SharedReg1110_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1110_out;
SharedReg617_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_57_cast <= SharedReg617_out;
SharedReg1118_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1118_out;
SharedReg1112_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1112_out;
SharedReg1157_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1157_out;
SharedReg1026_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1026_out;
SharedReg625_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_62_cast <= SharedReg625_out;
SharedReg622_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_63_cast <= SharedReg622_out;
SharedReg1078_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1078_out;
   MUX_Product32_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg95_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1165_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg617_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg617_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1129_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1144_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1130_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1131_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1146_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg618_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg618_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1134_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg913_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1149_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1055_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1056_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg88_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg931_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1170_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg88_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1005_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1059_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg935_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1139_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg265_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1109_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1009_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1169_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1167_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg269_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg94_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1012_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1065_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1122_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1126_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1014_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg272_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1016_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1068_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1069_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg628_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1097_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1098_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg944_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1100_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1127_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg940_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1053_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1102_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1162_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1116_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1110_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg617_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1118_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1112_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1157_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg622_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1026_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg625_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg622_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1078_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1141_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1128_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1054_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product32_2_impl_0_out);

   Delay1No104_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_2_impl_0_out,
                 Y => Delay1No104_out);

SharedReg1079_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1079_out;
SharedReg624_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg624_out;
SharedReg1138_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1138_out;
SharedReg625_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg625_out;
SharedReg626_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg626_out;
SharedReg621_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg621_out;
SharedReg1140_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1140_out;
SharedReg911_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg911_out;
SharedReg912_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg912_out;
SharedReg279_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg279_out;
SharedReg1142_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1142_out;
SharedReg1143_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1143_out;
SharedReg618_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg618_out;
SharedReg618_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg618_out;
SharedReg619_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg619_out;
SharedReg622_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg622_out;
SharedReg618_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg618_out;
SharedReg1147_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg1147_out;
SharedReg1148_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1148_out;
SharedReg619_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg619_out;
SharedReg619_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg619_out;
SharedReg953_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg953_out;
SharedReg950_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg950_out;
SharedReg1095_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1095_out;
SharedReg1057_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1057_out;
SharedReg931_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg931_out;
SharedReg1058_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1058_out;
SharedReg260_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg260_out;
SharedReg89_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_29_cast <= SharedReg89_out;
SharedReg1171_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_30_cast <= SharedReg1171_out;
SharedReg1060_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_31_cast <= SharedReg1060_out;
SharedReg621_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_32_cast <= SharedReg621_out;
SharedReg939_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_33_cast <= SharedReg939_out;
SharedReg934_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_34_cast <= SharedReg934_out;
SharedReg935_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_35_cast <= SharedReg935_out;
SharedReg1063_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_36_cast <= SharedReg1063_out;
SharedReg1064_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_37_cast <= SharedReg1064_out;
SharedReg630_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_38_cast <= SharedReg630_out;
SharedReg97_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_39_cast <= SharedReg97_out;
SharedReg628_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_40_cast <= SharedReg628_out;
SharedReg274_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_41_cast <= SharedReg274_out;
SharedReg1066_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_42_cast <= SharedReg1066_out;
SharedReg99_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_43_cast <= SharedReg99_out;
SharedReg275_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_44_cast <= SharedReg275_out;
SharedReg100_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_45_cast <= SharedReg100_out;
SharedReg1096_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_46_cast <= SharedReg1096_out;
SharedReg98_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_47_cast <= SharedReg98_out;
SharedReg629_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_48_cast <= SharedReg629_out;
SharedReg1099_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_49_cast <= SharedReg1099_out;
SharedReg944_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_50_cast <= SharedReg944_out;
SharedReg1101_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_51_cast <= SharedReg1101_out;
SharedReg941_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_52_cast <= SharedReg941_out;
SharedReg269_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_53_cast <= SharedReg269_out;
SharedReg906_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_54_cast <= SharedReg906_out;
SharedReg906_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_55_cast <= SharedReg906_out;
SharedReg907_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_56_cast <= SharedReg907_out;
SharedReg1163_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1163_out;
SharedReg931_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_58_cast <= SharedReg931_out;
SharedReg932_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_59_cast <= SharedReg932_out;
SharedReg620_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_60_cast <= SharedReg620_out;
SharedReg91_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_61_cast <= SharedReg91_out;
SharedReg1164_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_62_cast <= SharedReg1164_out;
SharedReg1077_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_63_cast <= SharedReg1077_out;
SharedReg938_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_64_cast <= SharedReg938_out;
   MUX_Product32_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1079_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg624_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1142_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1143_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg618_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg618_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg619_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg622_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg618_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1147_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1148_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg619_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1138_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg619_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg953_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg950_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1095_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1057_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg931_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1058_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg260_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg89_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1171_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg625_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1060_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg621_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg939_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg934_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg935_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1063_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1064_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg630_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg97_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg628_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg626_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg274_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1066_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg99_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg275_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg100_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1096_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg98_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg629_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1099_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg944_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg621_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1101_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg941_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg269_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg906_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg906_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg907_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1163_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg931_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg932_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg620_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1140_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg91_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1164_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1077_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg938_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg911_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg912_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg279_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product32_2_impl_1_out);

   Delay1No105_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_2_impl_1_out,
                 Y => Delay1No105_out);

Delay1No106_out_to_Product32_3_impl_parent_implementedSystem_port_0_cast <= Delay1No106_out;
Delay1No107_out_to_Product32_3_impl_parent_implementedSystem_port_1_cast <= Delay1No107_out;
   Product32_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_3_impl_out,
                 X => Delay1No106_out_to_Product32_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No107_out_to_Product32_3_impl_parent_implementedSystem_port_1_cast);

SharedReg1110_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1110_out;
SharedReg931_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg931_out;
SharedReg1118_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1118_out;
SharedReg1112_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1112_out;
SharedReg1157_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1157_out;
SharedReg1026_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1026_out;
SharedReg939_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg939_out;
SharedReg936_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg936_out;
SharedReg1078_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1078_out;
SharedReg268_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg268_out;
SharedReg1165_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1165_out;
SharedReg624_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg624_out;
SharedReg1139_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1139_out;
SharedReg1126_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1126_out;
SharedReg1127_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1127_out;
SharedReg645_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg645_out;
SharedReg1141_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1141_out;
SharedReg1128_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1128_out;
SharedReg1054_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1054_out;
SharedReg640_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg640_out;
SharedReg640_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg640_out;
SharedReg1129_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1129_out;
SharedReg1144_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1144_out;
SharedReg1130_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1130_out;
SharedReg1131_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1131_out;
SharedReg1146_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1146_out;
SharedReg641_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg641_out;
SharedReg641_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg641_out;
SharedReg1134_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1134_out;
SharedReg1149_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_30_cast <= SharedReg1149_out;
SharedReg1055_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1055_out;
SharedReg1056_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1056_out;
SharedReg260_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_33_cast <= SharedReg260_out;
SharedReg855_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_34_cast <= SharedReg855_out;
SharedReg1170_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1170_out;
SharedReg114_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_36_cast <= SharedReg114_out;
SharedReg1005_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1005_out;
SharedReg1059_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1059_out;
SharedReg859_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_39_cast <= SharedReg859_out;
SharedReg290_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_40_cast <= SharedReg290_out;
SharedReg1109_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1109_out;
SharedReg1009_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1009_out;
SharedReg1169_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1169_out;
SharedReg1167_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1167_out;
SharedReg294_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_45_cast <= SharedReg294_out;
SharedReg120_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_46_cast <= SharedReg120_out;
SharedReg1012_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1012_out;
SharedReg1065_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1065_out;
SharedReg1122_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1122_out;
SharedReg1014_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1014_out;
SharedReg297_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_51_cast <= SharedReg297_out;
SharedReg1016_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1016_out;
SharedReg1068_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1068_out;
SharedReg1069_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1069_out;
SharedReg650_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_55_cast <= SharedReg650_out;
SharedReg1097_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1097_out;
SharedReg1098_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1098_out;
SharedReg869_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_58_cast <= SharedReg869_out;
SharedReg1100_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1100_out;
SharedReg864_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_60_cast <= SharedReg864_out;
SharedReg1053_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1053_out;
SharedReg1102_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1102_out;
SharedReg1162_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1162_out;
SharedReg1116_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_64_cast <= SharedReg1116_out;
   MUX_Product32_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1110_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg931_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1165_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg624_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1139_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1126_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1127_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg645_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1141_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1128_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1054_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg640_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1118_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg640_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1129_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1144_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1130_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1131_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1146_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg641_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg641_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1134_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1149_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1112_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1055_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1056_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg260_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg855_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1170_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg114_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1005_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1059_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg859_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg290_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1157_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1109_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1009_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1169_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1167_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg294_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg120_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1012_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1065_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1122_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1014_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1026_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg297_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1016_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1068_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1069_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg650_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1097_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1098_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg869_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1100_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg864_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg939_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1053_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1102_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1162_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1116_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg936_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1078_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg268_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product32_3_impl_0_out);

   Delay1No106_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_3_impl_0_out,
                 Y => Delay1No106_out);

SharedReg618_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg618_out;
SharedReg1163_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1163_out;
SharedReg640_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg640_out;
SharedReg641_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg641_out;
SharedReg934_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg934_out;
SharedReg264_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg264_out;
SharedReg1164_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1164_out;
SharedReg1077_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1077_out;
SharedReg647_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg647_out;
SharedReg1079_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1079_out;
SharedReg938_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg938_out;
SharedReg1138_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1138_out;
SharedReg939_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg939_out;
SharedReg940_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg940_out;
SharedReg644_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg644_out;
SharedReg1140_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1140_out;
SharedReg936_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg936_out;
SharedReg937_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg937_out;
SharedReg305_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg305_out;
SharedReg1142_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1142_out;
SharedReg1143_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1143_out;
SharedReg641_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg641_out;
SharedReg641_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg641_out;
SharedReg642_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg642_out;
SharedReg645_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg645_out;
SharedReg641_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg641_out;
SharedReg1147_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg1147_out;
SharedReg1148_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1148_out;
SharedReg642_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_29_cast <= SharedReg642_out;
SharedReg642_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_30_cast <= SharedReg642_out;
SharedReg878_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_31_cast <= SharedReg878_out;
SharedReg875_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_32_cast <= SharedReg875_out;
SharedReg1095_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_33_cast <= SharedReg1095_out;
SharedReg1057_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_34_cast <= SharedReg1057_out;
SharedReg855_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_35_cast <= SharedReg855_out;
SharedReg1058_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_36_cast <= SharedReg1058_out;
SharedReg285_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_37_cast <= SharedReg285_out;
SharedReg115_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_38_cast <= SharedReg115_out;
SharedReg1171_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_39_cast <= SharedReg1171_out;
SharedReg1060_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_40_cast <= SharedReg1060_out;
SharedReg644_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_41_cast <= SharedReg644_out;
SharedReg863_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_42_cast <= SharedReg863_out;
SharedReg858_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_43_cast <= SharedReg858_out;
SharedReg859_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_44_cast <= SharedReg859_out;
SharedReg1063_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_45_cast <= SharedReg1063_out;
SharedReg1064_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_46_cast <= SharedReg1064_out;
SharedReg651_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_47_cast <= SharedReg651_out;
SharedReg123_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_48_cast <= SharedReg123_out;
SharedReg650_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_49_cast <= SharedReg650_out;
SharedReg299_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_50_cast <= SharedReg299_out;
SharedReg1066_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_51_cast <= SharedReg1066_out;
SharedReg124_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_52_cast <= SharedReg124_out;
SharedReg300_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_53_cast <= SharedReg300_out;
SharedReg125_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_54_cast <= SharedReg125_out;
SharedReg1096_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_55_cast <= SharedReg1096_out;
SharedReg271_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_56_cast <= SharedReg271_out;
SharedReg943_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_57_cast <= SharedReg943_out;
SharedReg1099_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_58_cast <= SharedReg1099_out;
SharedReg652_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_59_cast <= SharedReg652_out;
SharedReg1101_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_60_cast <= SharedReg1101_out;
SharedReg865_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_61_cast <= SharedReg865_out;
SharedReg294_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_62_cast <= SharedReg294_out;
SharedReg617_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_63_cast <= SharedReg617_out;
SharedReg617_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_64_cast <= SharedReg617_out;
   MUX_Product32_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg618_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1163_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg938_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1138_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg939_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg940_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg644_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1140_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg936_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg937_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg305_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1142_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg640_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1143_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg641_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg641_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg642_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg645_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg641_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1147_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1148_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg642_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg642_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg641_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg878_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg875_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1095_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1057_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg855_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1058_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg285_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg115_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1171_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1060_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg934_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg644_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg863_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg858_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg859_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1063_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1064_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg651_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg123_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg650_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg299_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg264_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1066_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg124_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg300_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg125_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1096_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg271_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg943_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1099_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg652_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1101_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1164_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg865_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg294_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg617_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg617_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1077_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg647_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1079_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product32_3_impl_1_out);

   Delay1No107_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_3_impl_1_out,
                 Y => Delay1No107_out);

Delay1No108_out_to_Product32_4_impl_parent_implementedSystem_port_0_cast <= Delay1No108_out;
Delay1No109_out_to_Product32_4_impl_parent_implementedSystem_port_1_cast <= Delay1No109_out;
   Product32_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_4_impl_out,
                 X => Delay1No108_out_to_Product32_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No109_out_to_Product32_4_impl_parent_implementedSystem_port_1_cast);

SharedReg1097_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1097_out;
SharedReg1098_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1098_out;
SharedReg698_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg698_out;
SharedReg1100_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1100_out;
SharedReg670_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg670_out;
SharedReg1053_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1053_out;
SharedReg1102_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1102_out;
SharedReg1162_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1162_out;
SharedReg1116_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1116_out;
SharedReg1110_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1110_out;
SharedReg855_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg855_out;
SharedReg1118_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1118_out;
SharedReg1112_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1112_out;
SharedReg1157_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1157_out;
SharedReg1026_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1026_out;
SharedReg863_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg863_out;
SharedReg860_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg860_out;
SharedReg1078_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1078_out;
SharedReg293_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg293_out;
SharedReg1165_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1165_out;
SharedReg647_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg647_out;
SharedReg1139_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1139_out;
SharedReg1126_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1126_out;
SharedReg1127_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1127_out;
SharedReg666_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg666_out;
SharedReg1141_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1141_out;
SharedReg1128_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1128_out;
SharedReg1054_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1054_out;
SharedReg661_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_29_cast <= SharedReg661_out;
SharedReg661_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_30_cast <= SharedReg661_out;
SharedReg1129_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1129_out;
SharedReg1144_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1144_out;
SharedReg1130_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1130_out;
SharedReg1131_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1131_out;
SharedReg1146_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1146_out;
SharedReg662_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_36_cast <= SharedReg662_out;
SharedReg662_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_37_cast <= SharedReg662_out;
SharedReg1134_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_38_cast <= SharedReg1134_out;
SharedReg1149_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1149_out;
SharedReg1055_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1055_out;
SharedReg1056_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1056_out;
SharedReg285_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_42_cast <= SharedReg285_out;
SharedReg685_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_43_cast <= SharedReg685_out;
SharedReg1170_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1170_out;
SharedReg285_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_45_cast <= SharedReg285_out;
SharedReg1005_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1005_out;
SharedReg1059_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1059_out;
SharedReg689_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_48_cast <= SharedReg689_out;
SharedReg315_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_49_cast <= SharedReg315_out;
SharedReg1109_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1109_out;
SharedReg1009_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1009_out;
SharedReg1169_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1169_out;
SharedReg1167_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1167_out;
SharedReg146_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_54_cast <= SharedReg146_out;
SharedReg144_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_55_cast <= SharedReg144_out;
SharedReg1012_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1012_out;
SharedReg1065_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1065_out;
SharedReg1122_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1122_out;
SharedReg1014_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1014_out;
SharedReg320_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_60_cast <= SharedReg320_out;
SharedReg1016_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1016_out;
SharedReg1068_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1068_out;
SharedReg1069_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1069_out;
SharedReg672_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_64_cast <= SharedReg672_out;
   MUX_Product32_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1097_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1098_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg855_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1118_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1112_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1157_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1026_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg863_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg860_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1078_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg293_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1165_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg698_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg647_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1139_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1126_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1127_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg666_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1141_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1128_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1054_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg661_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg661_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1100_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1129_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1144_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1130_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1131_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1146_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg662_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg662_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1134_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1149_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1055_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg670_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1056_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg285_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg685_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1170_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg285_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1005_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1059_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg689_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg315_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1109_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1053_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1009_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1169_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1167_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg146_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg144_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1012_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1065_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1122_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1014_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg320_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1102_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1016_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1068_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1069_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg672_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1162_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1116_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1110_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product32_4_impl_0_out);

   Delay1No108_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_4_impl_0_out,
                 Y => Delay1No108_out);

SharedReg296_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg296_out;
SharedReg867_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg867_out;
SharedReg1099_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1099_out;
SharedReg675_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg675_out;
SharedReg1101_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1101_out;
SharedReg671_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg671_out;
SharedReg146_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg146_out;
SharedReg640_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg640_out;
SharedReg640_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg640_out;
SharedReg641_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg641_out;
SharedReg1163_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1163_out;
SharedReg661_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg661_out;
SharedReg662_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg662_out;
SharedReg858_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg858_out;
SharedReg289_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg289_out;
SharedReg1164_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg1164_out;
SharedReg1077_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg1077_out;
SharedReg668_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg668_out;
SharedReg1079_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1079_out;
SharedReg862_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg862_out;
SharedReg1138_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg1138_out;
SharedReg863_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg863_out;
SharedReg864_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg864_out;
SharedReg665_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg665_out;
SharedReg1140_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1140_out;
SharedReg860_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg860_out;
SharedReg861_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg861_out;
SharedReg153_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg153_out;
SharedReg1142_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_29_cast <= SharedReg1142_out;
SharedReg1143_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_30_cast <= SharedReg1143_out;
SharedReg662_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_31_cast <= SharedReg662_out;
SharedReg662_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_32_cast <= SharedReg662_out;
SharedReg663_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_33_cast <= SharedReg663_out;
SharedReg666_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_34_cast <= SharedReg666_out;
SharedReg662_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_35_cast <= SharedReg662_out;
SharedReg1147_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_36_cast <= SharedReg1147_out;
SharedReg1148_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_37_cast <= SharedReg1148_out;
SharedReg663_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_38_cast <= SharedReg663_out;
SharedReg663_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_39_cast <= SharedReg663_out;
SharedReg681_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_40_cast <= SharedReg681_out;
SharedReg678_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_41_cast <= SharedReg678_out;
SharedReg1095_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_42_cast <= SharedReg1095_out;
SharedReg1057_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_43_cast <= SharedReg1057_out;
SharedReg685_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_44_cast <= SharedReg685_out;
SharedReg1058_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_45_cast <= SharedReg1058_out;
SharedReg285_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_46_cast <= SharedReg285_out;
SharedReg115_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_47_cast <= SharedReg115_out;
SharedReg1171_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_48_cast <= SharedReg1171_out;
SharedReg1060_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_49_cast <= SharedReg1060_out;
SharedReg644_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_50_cast <= SharedReg644_out;
SharedReg693_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_51_cast <= SharedReg693_out;
SharedReg688_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_52_cast <= SharedReg688_out;
SharedReg689_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_53_cast <= SharedReg689_out;
SharedReg1063_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_54_cast <= SharedReg1063_out;
SharedReg1064_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_55_cast <= SharedReg1064_out;
SharedReg674_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_56_cast <= SharedReg674_out;
SharedReg295_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_57_cast <= SharedReg295_out;
SharedReg866_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_58_cast <= SharedReg866_out;
SharedReg151_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_59_cast <= SharedReg151_out;
SharedReg1066_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_60_cast <= SharedReg1066_out;
SharedReg149_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_61_cast <= SharedReg149_out;
SharedReg152_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_62_cast <= SharedReg152_out;
SharedReg150_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_63_cast <= SharedReg150_out;
SharedReg1096_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_64_cast <= SharedReg1096_out;
   MUX_Product32_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg296_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg867_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1163_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg661_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg662_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg858_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg289_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1164_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1077_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg668_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1079_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg862_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1099_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1138_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg863_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg864_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg665_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1140_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg860_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg861_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg153_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1142_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1143_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg675_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg662_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg662_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg663_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg666_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg662_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1147_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1148_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg663_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg663_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg681_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1101_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg678_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1095_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1057_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg685_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1058_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg285_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg115_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1171_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1060_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg644_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg671_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg693_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg688_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg689_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1063_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1064_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg674_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg295_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg866_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg151_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1066_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg146_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg149_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg152_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg150_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1096_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg640_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg640_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg641_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product32_4_impl_1_out);

   Delay1No109_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_4_impl_1_out,
                 Y => Delay1No109_out);

Delay1No110_out_to_Product32_5_impl_parent_implementedSystem_port_0_cast <= Delay1No110_out;
Delay1No111_out_to_Product32_5_impl_parent_implementedSystem_port_1_cast <= Delay1No111_out;
   Product32_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_5_impl_out,
                 X => Delay1No110_out_to_Product32_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No111_out_to_Product32_5_impl_parent_implementedSystem_port_1_cast);

SharedReg1012_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1012_out;
SharedReg1065_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1065_out;
SharedReg1122_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1122_out;
SharedReg1014_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1014_out;
SharedReg198_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg198_out;
SharedReg1016_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1016_out;
SharedReg1068_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1068_out;
SharedReg1069_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1069_out;
SharedReg696_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg696_out;
SharedReg1097_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1097_out;
SharedReg1098_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1098_out;
SharedReg719_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg719_out;
SharedReg1100_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1100_out;
SharedReg694_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_14_cast <= SharedReg694_out;
SharedReg1053_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_15_cast <= SharedReg1053_out;
SharedReg1102_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1102_out;
SharedReg1162_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1162_out;
SharedReg1116_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1116_out;
SharedReg1110_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_19_cast <= SharedReg1110_out;
SharedReg685_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_20_cast <= SharedReg685_out;
SharedReg1118_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1118_out;
SharedReg1112_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_22_cast <= SharedReg1112_out;
SharedReg1157_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1157_out;
SharedReg1026_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1026_out;
SharedReg693_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_25_cast <= SharedReg693_out;
SharedReg690_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_26_cast <= SharedReg690_out;
SharedReg1078_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1078_out;
SharedReg317_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_28_cast <= SharedReg317_out;
SharedReg1165_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1165_out;
SharedReg862_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_30_cast <= SharedReg862_out;
SharedReg1139_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1139_out;
SharedReg1126_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1126_out;
SharedReg1127_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1127_out;
SharedReg712_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_34_cast <= SharedReg712_out;
SharedReg1141_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1141_out;
SharedReg1128_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_36_cast <= SharedReg1128_out;
SharedReg1054_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1054_out;
SharedReg707_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_38_cast <= SharedReg707_out;
SharedReg707_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_39_cast <= SharedReg707_out;
SharedReg1129_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_40_cast <= SharedReg1129_out;
SharedReg1144_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1144_out;
SharedReg1130_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1130_out;
SharedReg1131_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1131_out;
SharedReg1146_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_44_cast <= SharedReg1146_out;
SharedReg708_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_45_cast <= SharedReg708_out;
SharedReg686_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_46_cast <= SharedReg686_out;
SharedReg1134_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1134_out;
SharedReg1149_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_48_cast <= SharedReg1149_out;
SharedReg1055_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_49_cast <= SharedReg1055_out;
SharedReg1056_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1056_out;
SharedReg310_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_51_cast <= SharedReg310_out;
SharedReg882_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_52_cast <= SharedReg882_out;
SharedReg1170_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1170_out;
SharedReg310_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_54_cast <= SharedReg310_out;
SharedReg1005_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_55_cast <= SharedReg1005_out;
SharedReg1059_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_56_cast <= SharedReg1059_out;
SharedReg886_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_57_cast <= SharedReg886_out;
SharedReg191_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_58_cast <= SharedReg191_out;
SharedReg1109_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1109_out;
SharedReg1009_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1009_out;
SharedReg1169_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_61_cast <= SharedReg1169_out;
SharedReg1167_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_62_cast <= SharedReg1167_out;
SharedReg172_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_63_cast <= SharedReg172_out;
SharedReg170_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_64_cast <= SharedReg170_out;
   MUX_Product32_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1012_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1065_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1098_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg719_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1100_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg694_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1053_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1102_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1162_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1116_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1110_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg685_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1122_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1118_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1112_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1157_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1026_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg693_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg690_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1078_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg317_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1165_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg862_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1014_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1139_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1126_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1127_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg712_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1141_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1128_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1054_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg707_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg707_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1129_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg198_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1144_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1130_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1131_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1146_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg708_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg686_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1134_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1149_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1055_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1056_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1016_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg310_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg882_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1170_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg310_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1005_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1059_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg886_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg191_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1109_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1009_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1068_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1169_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1167_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg172_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg170_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1069_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg696_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1097_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product32_5_impl_0_out);

   Delay1No110_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_5_impl_0_out,
                 Y => Delay1No110_out);

SharedReg718_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg718_out;
SharedReg147_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg147_out;
SharedReg672_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg672_out;
SharedReg176_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg176_out;
SharedReg1066_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1066_out;
SharedReg174_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg174_out;
SharedReg323_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg323_out;
SharedReg175_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg175_out;
SharedReg1096_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1096_out;
SharedReg148_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg148_out;
SharedReg673_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg673_out;
SharedReg1099_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1099_out;
SharedReg698_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg698_out;
SharedReg1101_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_14_cast <= SharedReg1101_out;
SharedReg695_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_15_cast <= SharedReg695_out;
SharedReg172_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_16_cast <= SharedReg172_out;
SharedReg661_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_17_cast <= SharedReg661_out;
SharedReg661_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_18_cast <= SharedReg661_out;
SharedReg662_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_19_cast <= SharedReg662_out;
SharedReg1163_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_20_cast <= SharedReg1163_out;
SharedReg707_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_21_cast <= SharedReg707_out;
SharedReg708_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_22_cast <= SharedReg708_out;
SharedReg688_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_23_cast <= SharedReg688_out;
SharedReg314_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_24_cast <= SharedReg314_out;
SharedReg1164_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_25_cast <= SharedReg1164_out;
SharedReg1077_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_26_cast <= SharedReg1077_out;
SharedReg714_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_27_cast <= SharedReg714_out;
SharedReg1079_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_28_cast <= SharedReg1079_out;
SharedReg692_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_29_cast <= SharedReg692_out;
SharedReg1138_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_30_cast <= SharedReg1138_out;
SharedReg669_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_31_cast <= SharedReg669_out;
SharedReg670_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_32_cast <= SharedReg670_out;
SharedReg711_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_33_cast <= SharedReg711_out;
SharedReg1140_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_34_cast <= SharedReg1140_out;
SharedReg690_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_35_cast <= SharedReg690_out;
SharedReg691_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_36_cast <= SharedReg691_out;
SharedReg178_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_37_cast <= SharedReg178_out;
SharedReg1142_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_38_cast <= SharedReg1142_out;
SharedReg1143_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_39_cast <= SharedReg1143_out;
SharedReg708_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_40_cast <= SharedReg708_out;
SharedReg708_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_41_cast <= SharedReg708_out;
SharedReg709_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_42_cast <= SharedReg709_out;
SharedReg712_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_43_cast <= SharedReg712_out;
SharedReg708_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_44_cast <= SharedReg708_out;
SharedReg1147_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_45_cast <= SharedReg1147_out;
SharedReg1148_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_46_cast <= SharedReg1148_out;
SharedReg687_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_47_cast <= SharedReg687_out;
SharedReg663_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_48_cast <= SharedReg663_out;
SharedReg725_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_49_cast <= SharedReg725_out;
SharedReg722_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_50_cast <= SharedReg722_out;
SharedReg1095_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_51_cast <= SharedReg1095_out;
SharedReg1057_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_52_cast <= SharedReg1057_out;
SharedReg882_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_53_cast <= SharedReg882_out;
SharedReg1058_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_54_cast <= SharedReg1058_out;
SharedReg310_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_55_cast <= SharedReg310_out;
SharedReg140_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_56_cast <= SharedReg140_out;
SharedReg1171_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_57_cast <= SharedReg1171_out;
SharedReg1060_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_58_cast <= SharedReg1060_out;
SharedReg665_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_59_cast <= SharedReg665_out;
SharedReg890_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_60_cast <= SharedReg890_out;
SharedReg885_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_61_cast <= SharedReg885_out;
SharedReg886_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_62_cast <= SharedReg886_out;
SharedReg1063_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_63_cast <= SharedReg1063_out;
SharedReg1064_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_64_cast <= SharedReg1064_out;
   MUX_Product32_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg718_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg147_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg673_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1099_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg698_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1101_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg695_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg172_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg661_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg661_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg662_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1163_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg672_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg707_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg708_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg688_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg314_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1164_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1077_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg714_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1079_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg692_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1138_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg176_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg669_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg670_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg711_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1140_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg690_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg691_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg178_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1142_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1143_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg708_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1066_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg708_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg709_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg712_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg708_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1147_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1148_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg687_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg663_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg725_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg722_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg174_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1095_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1057_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg882_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1058_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg310_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg140_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1171_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1060_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg665_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg890_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg323_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg885_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg886_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1063_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1064_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg175_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1096_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg148_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product32_5_impl_1_out);

   Delay1No111_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_5_impl_1_out,
                 Y => Delay1No111_out);

Delay1No112_out_to_Product32_6_impl_parent_implementedSystem_port_0_cast <= Delay1No112_out;
Delay1No113_out_to_Product32_6_impl_parent_implementedSystem_port_1_cast <= Delay1No113_out;
   Product32_6_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_6_impl_out,
                 X => Delay1No112_out_to_Product32_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No113_out_to_Product32_6_impl_parent_implementedSystem_port_1_cast);

SharedReg1005_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1005_out;
SharedReg1059_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1059_out;
SharedReg886_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg886_out;
SharedReg191_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg191_out;
SharedReg1109_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1109_out;
SharedReg1009_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1009_out;
SharedReg1169_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1169_out;
SharedReg1167_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1167_out;
SharedReg172_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg172_out;
SharedReg193_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg193_out;
SharedReg1012_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1012_out;
SharedReg1065_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1065_out;
SharedReg1122_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1122_out;
SharedReg1014_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_14_cast <= SharedReg1014_out;
SharedReg342_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_15_cast <= SharedReg342_out;
SharedReg1016_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1016_out;
SharedReg1068_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_17_cast <= SharedReg1068_out;
SharedReg1069_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_18_cast <= SharedReg1069_out;
SharedReg717_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_19_cast <= SharedReg717_out;
SharedReg1097_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1097_out;
SharedReg1098_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_21_cast <= SharedReg1098_out;
SharedReg895_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_22_cast <= SharedReg895_out;
SharedReg1100_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_23_cast <= SharedReg1100_out;
SharedReg992_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_24_cast <= SharedReg992_out;
SharedReg1053_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_25_cast <= SharedReg1053_out;
SharedReg1102_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_26_cast <= SharedReg1102_out;
SharedReg1162_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_27_cast <= SharedReg1162_out;
SharedReg1116_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_28_cast <= SharedReg1116_out;
SharedReg1110_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1110_out;
SharedReg882_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_30_cast <= SharedReg882_out;
SharedReg1118_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_31_cast <= SharedReg1118_out;
SharedReg1112_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_32_cast <= SharedReg1112_out;
SharedReg1157_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_33_cast <= SharedReg1157_out;
SharedReg1026_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_34_cast <= SharedReg1026_out;
SharedReg715_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_35_cast <= SharedReg715_out;
SharedReg887_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_36_cast <= SharedReg887_out;
SharedReg1078_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_37_cast <= SharedReg1078_out;
SharedReg194_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_38_cast <= SharedReg194_out;
SharedReg1165_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_39_cast <= SharedReg1165_out;
SharedReg889_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_40_cast <= SharedReg889_out;
SharedReg1139_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_41_cast <= SharedReg1139_out;
SharedReg1126_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_42_cast <= SharedReg1126_out;
SharedReg1127_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_43_cast <= SharedReg1127_out;
SharedReg988_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_44_cast <= SharedReg988_out;
SharedReg1141_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_45_cast <= SharedReg1141_out;
SharedReg1128_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_46_cast <= SharedReg1128_out;
SharedReg1054_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1054_out;
SharedReg983_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_48_cast <= SharedReg983_out;
SharedReg983_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_49_cast <= SharedReg983_out;
SharedReg1129_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_50_cast <= SharedReg1129_out;
SharedReg1144_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_51_cast <= SharedReg1144_out;
SharedReg1130_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_52_cast <= SharedReg1130_out;
SharedReg1131_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_53_cast <= SharedReg1131_out;
SharedReg1146_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_54_cast <= SharedReg1146_out;
SharedReg883_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_55_cast <= SharedReg883_out;
SharedReg708_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_56_cast <= SharedReg708_out;
SharedReg1134_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_57_cast <= SharedReg1134_out;
SharedReg1149_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_58_cast <= SharedReg1149_out;
SharedReg1055_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_59_cast <= SharedReg1055_out;
SharedReg1056_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_60_cast <= SharedReg1056_out;
SharedReg186_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_61_cast <= SharedReg186_out;
SharedReg983_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_62_cast <= SharedReg983_out;
SharedReg1170_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_63_cast <= SharedReg1170_out;
SharedReg310_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_64_cast <= SharedReg310_out;
   MUX_Product32_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1005_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1059_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1012_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1065_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1122_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg1014_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg342_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1016_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg1068_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg1069_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg717_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1097_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg886_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg1098_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg895_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg1100_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg992_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg1053_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg1102_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg1162_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg1116_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1110_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg882_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg191_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg1118_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg1112_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg1157_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg1026_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg715_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg887_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg1078_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg194_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg1165_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg889_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg1109_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1139_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg1126_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg1127_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg988_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg1141_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg1128_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1054_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg983_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg983_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg1129_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg1009_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg1144_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg1130_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg1131_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg1146_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg883_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg708_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg1134_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg1149_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg1055_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg1056_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg1169_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg186_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg983_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg1170_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg310_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg1167_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg172_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg193_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product32_6_impl_0_out);

   Delay1No112_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_6_impl_0_out,
                 Y => Delay1No112_out);

SharedReg163_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg163_out;
SharedReg311_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg311_out;
SharedReg1171_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1171_out;
SharedReg1060_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1060_out;
SharedReg689_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg689_out;
SharedReg991_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg991_out;
SharedReg885_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg885_out;
SharedReg886_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg886_out;
SharedReg1063_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1063_out;
SharedReg1064_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1064_out;
SharedReg894_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg894_out;
SharedReg196_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg196_out;
SharedReg892_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_13_cast <= SharedReg892_out;
SharedReg176_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_14_cast <= SharedReg176_out;
SharedReg1066_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_15_cast <= SharedReg1066_out;
SharedReg198_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_16_cast <= SharedReg198_out;
SharedReg343_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_17_cast <= SharedReg343_out;
SharedReg321_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_18_cast <= SharedReg321_out;
SharedReg1096_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_19_cast <= SharedReg1096_out;
SharedReg319_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_20_cast <= SharedReg319_out;
SharedReg697_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_21_cast <= SharedReg697_out;
SharedReg1099_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_22_cast <= SharedReg1099_out;
SharedReg719_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_23_cast <= SharedReg719_out;
SharedReg1101_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_24_cast <= SharedReg1101_out;
SharedReg993_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_25_cast <= SharedReg993_out;
SharedReg195_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_26_cast <= SharedReg195_out;
SharedReg685_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_27_cast <= SharedReg685_out;
SharedReg707_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_28_cast <= SharedReg707_out;
SharedReg708_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_29_cast <= SharedReg708_out;
SharedReg1163_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_30_cast <= SharedReg1163_out;
SharedReg983_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_31_cast <= SharedReg983_out;
SharedReg984_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_32_cast <= SharedReg984_out;
SharedReg885_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_33_cast <= SharedReg885_out;
SharedReg190_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_34_cast <= SharedReg190_out;
SharedReg1164_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_35_cast <= SharedReg1164_out;
SharedReg1077_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_36_cast <= SharedReg1077_out;
SharedReg990_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_37_cast <= SharedReg990_out;
SharedReg1079_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_38_cast <= SharedReg1079_out;
SharedReg692_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_39_cast <= SharedReg692_out;
SharedReg1138_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_40_cast <= SharedReg1138_out;
SharedReg991_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_41_cast <= SharedReg991_out;
SharedReg992_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_42_cast <= SharedReg992_out;
SharedReg987_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_43_cast <= SharedReg987_out;
SharedReg1140_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_44_cast <= SharedReg1140_out;
SharedReg887_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_45_cast <= SharedReg887_out;
SharedReg888_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_46_cast <= SharedReg888_out;
SharedReg204_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_47_cast <= SharedReg204_out;
SharedReg1142_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_48_cast <= SharedReg1142_out;
SharedReg1143_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_49_cast <= SharedReg1143_out;
SharedReg984_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_50_cast <= SharedReg984_out;
SharedReg883_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_51_cast <= SharedReg883_out;
SharedReg884_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_52_cast <= SharedReg884_out;
SharedReg988_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_53_cast <= SharedReg988_out;
SharedReg984_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_54_cast <= SharedReg984_out;
SharedReg1147_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_55_cast <= SharedReg1147_out;
SharedReg1148_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_56_cast <= SharedReg1148_out;
SharedReg709_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_57_cast <= SharedReg709_out;
SharedReg709_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_58_cast <= SharedReg709_out;
SharedReg902_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_59_cast <= SharedReg902_out;
SharedReg998_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_60_cast <= SharedReg998_out;
SharedReg1095_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_61_cast <= SharedReg1095_out;
SharedReg1057_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_62_cast <= SharedReg1057_out;
SharedReg882_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_63_cast <= SharedReg882_out;
SharedReg1058_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_64_cast <= SharedReg1058_out;
   MUX_Product32_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg163_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg311_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg894_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg196_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg892_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg176_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg1066_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg198_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg343_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg321_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg1096_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg319_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg1171_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg697_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg1099_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg719_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1101_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg993_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg195_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg685_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg707_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg708_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg1163_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg1060_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg983_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg984_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg885_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg190_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1164_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg1077_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg990_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg1079_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg692_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg1138_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg689_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg991_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg992_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg987_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg1140_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg887_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg888_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg204_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg1142_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg1143_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg984_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg991_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg883_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg884_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg988_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg984_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg1147_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg1148_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg709_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg709_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg902_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg998_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg885_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg1095_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg1057_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg882_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg1058_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg886_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1063_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1064_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Product32_6_impl_1_out);

   Delay1No113_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_6_impl_1_out,
                 Y => Delay1No113_out);

Delay1No114_out_to_Subtract3_4_impl_parent_implementedSystem_port_0_cast <= Delay1No114_out;
Delay1No115_out_to_Subtract3_4_impl_parent_implementedSystem_port_1_cast <= Delay1No115_out;
   Subtract3_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract3_4_impl_out,
                 X => Delay1No114_out_to_Subtract3_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No115_out_to_Subtract3_4_impl_parent_implementedSystem_port_1_cast);

SharedReg522_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg522_out;
SharedReg519_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg519_out;
SharedReg139_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg139_out;
SharedReg312_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg312_out;
SharedReg426_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg426_out;
SharedReg139_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg139_out;
SharedReg149_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg149_out;
SharedReg857_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg857_out;
SharedReg868_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg868_out;
SharedReg414_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg414_out;
SharedReg523_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg523_out;
SharedReg522_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg522_out;
SharedReg425_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg425_out;
SharedReg665_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg665_out;
SharedReg802_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg802_out;
SharedReg655_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg655_out;
SharedReg411_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg411_out;
SharedReg302_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg302_out;
SharedReg288_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg288_out;
SharedReg410_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg410_out;
SharedReg142_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg142_out;
SharedReg410_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg410_out;
SharedReg412_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg412_out;
SharedReg519_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg519_out;
SharedReg646_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg646_out;
SharedReg412_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg412_out;
SharedReg820_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg820_out;
SharedReg783_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg783_out;
SharedReg1_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_29_cast <= SharedReg1_out;
SharedReg3_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_30_cast <= SharedReg3_out;
SharedReg17_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_31_cast <= SharedReg17_out;
SharedReg6_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_32_cast <= SharedReg6_out;
SharedReg11_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_33_cast <= SharedReg11_out;
SharedReg12_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_34_cast <= SharedReg12_out;
SharedReg16_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_35_cast <= SharedReg16_out;
SharedReg410_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_36_cast <= SharedReg410_out;
SharedReg509_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_37_cast <= SharedReg509_out;
SharedReg506_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_38_cast <= SharedReg506_out;
SharedReg122_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_39_cast <= SharedReg122_out;
SharedReg14_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_40_cast <= SharedReg14_out;
SharedReg6_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_41_cast <= SharedReg6_out;
SharedReg7_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_42_cast <= SharedReg7_out;
SharedReg506_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_43_cast <= SharedReg506_out;
SharedReg404_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_44_cast <= SharedReg404_out;
SharedReg8_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_45_cast <= SharedReg8_out;
SharedReg278_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_46_cast <= SharedReg278_out;
SharedReg948_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_47_cast <= SharedReg948_out;
SharedReg948_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_48_cast <= SharedReg948_out;
SharedReg654_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_49_cast <= SharedReg654_out;
SharedReg813_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_50_cast <= SharedReg813_out;
SharedReg422_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_51_cast <= SharedReg422_out;
SharedReg134_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_52_cast <= SharedReg134_out;
SharedReg644_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_53_cast <= SharedReg644_out;
SharedReg503_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_54_cast <= SharedReg503_out;
SharedReg802_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_55_cast <= SharedReg802_out;
SharedReg410_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_56_cast <= SharedReg410_out;
SharedReg801_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_57_cast <= SharedReg801_out;
SharedReg287_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_58_cast <= SharedReg287_out;
SharedReg547_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_59_cast <= SharedReg547_out;
SharedReg535_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_60_cast <= SharedReg535_out;
SharedReg313_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_61_cast <= SharedReg313_out;
SharedReg410_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_62_cast <= SharedReg410_out;
SharedReg416_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_63_cast <= SharedReg416_out;
SharedReg315_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_64_cast <= SharedReg315_out;
   MUX_Subtract3_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg522_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg519_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg523_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg522_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg425_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg665_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg802_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg655_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg411_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg302_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg288_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg410_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg139_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg142_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg410_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg412_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg519_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg646_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg412_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg820_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg783_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg1_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg3_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg312_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg17_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg6_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg11_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg12_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg16_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg410_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg509_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg506_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg122_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg14_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg426_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg6_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg7_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg506_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg404_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg8_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg278_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg948_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg948_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg654_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg813_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg139_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg422_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg134_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg644_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg503_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg802_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg410_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg801_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg287_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg547_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg535_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg149_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg313_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg410_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg416_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg315_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg857_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg868_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg414_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract3_4_impl_0_out);

   Delay1No114_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_4_impl_0_out,
                 Y => Delay1No114_out);

SharedReg519_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg519_out;
SharedReg803_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg803_out;
SharedReg143_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg143_out;
SharedReg184_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg184_out;
SharedReg535_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg535_out;
SharedReg141_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg141_out;
SharedReg285_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg285_out;
SharedReg665_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg665_out;
SharedReg931_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg931_out;
SharedReg817_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg817_out;
SharedReg808_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg808_out;
SharedReg806_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg806_out;
SharedReg435_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg435_out;
SharedReg859_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg859_out;
SharedReg519_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg519_out;
SharedReg662_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg662_out;
SharedReg519_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg519_out;
SharedReg139_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg139_out;
SharedReg155_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg155_out;
SharedReg520_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg520_out;
SharedReg160_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg160_out;
SharedReg802_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg802_out;
SharedReg519_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg519_out;
SharedReg810_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg810_out;
SharedReg855_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg855_out;
SharedReg804_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg804_out;
SharedReg535_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg535_out;
SharedReg786_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg786_out;
SharedReg19_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_29_cast <= SharedReg19_out;
SharedReg21_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_30_cast <= SharedReg21_out;
SharedReg35_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_31_cast <= SharedReg35_out;
SharedReg24_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_32_cast <= SharedReg24_out;
SharedReg29_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_33_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_34_cast <= SharedReg30_out;
SharedReg34_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_35_cast <= SharedReg34_out;
SharedReg521_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_36_cast <= SharedReg521_out;
SharedReg789_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_37_cast <= SharedReg789_out;
SharedReg789_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_38_cast <= SharedReg789_out;
SharedReg123_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_39_cast <= SharedReg123_out;
SharedReg32_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_40_cast <= SharedReg32_out;
SharedReg24_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_41_cast <= SharedReg24_out;
SharedReg25_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_42_cast <= SharedReg25_out;
SharedReg783_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_43_cast <= SharedReg783_out;
SharedReg402_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_44_cast <= SharedReg402_out;
SharedReg26_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_45_cast <= SharedReg26_out;
SharedReg88_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_46_cast <= SharedReg88_out;
SharedReg932_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_47_cast <= SharedReg932_out;
SharedReg619_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_48_cast <= SharedReg619_out;
SharedReg676_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_49_cast <= SharedReg676_out;
SharedReg816_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_50_cast <= SharedReg816_out;
Delay43No11_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_51_cast <= Delay43No11_out;
SharedReg266_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_52_cast <= SharedReg266_out;
Delay76No3_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_53_cast <= Delay76No3_out;
SharedReg788_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_54_cast <= SharedReg788_out;
SharedReg410_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_55_cast <= SharedReg410_out;
SharedReg804_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_56_cast <= SharedReg804_out;
SharedReg418_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_57_cast <= SharedReg418_out;
SharedReg161_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_58_cast <= SharedReg161_out;
SharedReg437_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_59_cast <= SharedReg437_out;
SharedReg821_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_60_cast <= SharedReg821_out;
SharedReg308_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_61_cast <= SharedReg308_out;
SharedReg411_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_62_cast <= SharedReg411_out;
SharedReg410_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_63_cast <= SharedReg410_out;
Delay77No4_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_64_cast <= Delay77No4_out;
   MUX_Subtract3_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg519_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg803_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg808_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg806_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg435_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg859_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg519_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg662_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg519_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg139_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg155_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg520_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg143_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg160_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg802_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg519_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg810_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg855_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg804_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg535_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg786_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg19_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg21_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg184_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg35_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg24_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg29_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg30_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg34_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg521_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg789_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg789_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg123_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg32_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg535_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg24_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg25_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg783_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg402_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg26_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg88_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg932_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg619_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg676_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg816_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg141_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => Delay43No11_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg266_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => Delay76No3_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg788_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg410_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg804_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg418_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg161_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg437_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg821_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg285_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg308_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg411_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg410_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => Delay77No4_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg665_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg931_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg817_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract3_4_impl_1_out);

   Delay1No115_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_4_impl_1_out,
                 Y => Delay1No115_out);

Delay1No116_out_to_Subtract3_6_impl_parent_implementedSystem_port_0_cast <= Delay1No116_out;
Delay1No117_out_to_Subtract3_6_impl_parent_implementedSystem_port_1_cast <= Delay1No117_out;
   Subtract3_6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract3_6_impl_out,
                 X => Delay1No116_out_to_Subtract3_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No117_out_to_Subtract3_6_impl_parent_implementedSystem_port_1_cast);

SharedReg_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg_out;
SharedReg1_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1_out;
SharedReg3_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg3_out;
SharedReg3_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg3_out;
SharedReg7_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg7_out;
SharedReg10_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg10_out;
SharedReg12_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg12_out;
SharedReg13_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg13_out;
SharedReg16_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg16_out;
SharedReg16_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg16_out;
SharedReg320_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg320_out;
SharedReg721_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg721_out;
SharedReg440_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_13_cast <= SharedReg440_out;
SharedReg838_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_14_cast <= SharedReg838_out;
SharedReg440_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_15_cast <= SharedReg440_out;
SharedReg441_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_16_cast <= SharedReg441_out;
SharedReg441_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_17_cast <= SharedReg441_out;
SharedReg888_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_18_cast <= SharedReg888_out;
SharedReg202_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_19_cast <= SharedReg202_out;
SharedReg551_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_20_cast <= SharedReg551_out;
SharedReg897_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_21_cast <= SharedReg897_out;
SharedReg340_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_22_cast <= SharedReg340_out;
SharedReg440_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_23_cast <= SharedReg440_out;
SharedReg838_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_24_cast <= SharedReg838_out;
SharedReg888_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_25_cast <= SharedReg888_out;
SharedReg193_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_26_cast <= SharedReg193_out;
SharedReg838_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_27_cast <= SharedReg838_out;
SharedReg335_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_28_cast <= SharedReg335_out;
SharedReg851_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_29_cast <= SharedReg851_out;
SharedReg551_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_30_cast <= SharedReg551_out;
SharedReg332_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_31_cast <= SharedReg332_out;
SharedReg554_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_32_cast <= SharedReg554_out;
SharedReg445_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_33_cast <= SharedReg445_out;
SharedReg448_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_34_cast <= SharedReg448_out;
SharedReg989_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_35_cast <= SharedReg989_out;
SharedReg444_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_36_cast <= SharedReg444_out;
SharedReg440_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_37_cast <= SharedReg440_out;
SharedReg845_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_38_cast <= SharedReg845_out;
SharedReg189_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_39_cast <= SharedReg189_out;
SharedReg555_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_40_cast <= SharedReg555_out;
SharedReg440_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_41_cast <= SharedReg440_out;
SharedReg987_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_42_cast <= SharedReg987_out;
SharedReg440_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_43_cast <= SharedReg440_out;
SharedReg554_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_44_cast <= SharedReg554_out;
SharedReg886_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_45_cast <= SharedReg886_out;
SharedReg819_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_46_cast <= SharedReg819_out;
SharedReg338_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_47_cast <= SharedReg338_out;
   MUX_Subtract3_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_47_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg320_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg721_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg440_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg838_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg440_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg441_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg441_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg888_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg202_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg551_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg3_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg897_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg340_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg440_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg838_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg888_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg193_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg838_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg335_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg851_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg551_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg3_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg332_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg554_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg445_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg448_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg989_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg444_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg440_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg845_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg189_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg555_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg7_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg440_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg987_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg440_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg554_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg886_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg819_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg338_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_47_cast,
                 iS_5 => SharedReg10_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg12_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg13_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg16_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg16_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Subtract3_6_impl_0_LUT_out,
                 oMux => MUX_Subtract3_6_impl_0_out);

   Delay1No116_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_6_impl_0_out,
                 Y => Delay1No116_out);

SharedReg25_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg25_out;
SharedReg18_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg18_out;
SharedReg19_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg19_out;
SharedReg21_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg21_out;
SharedReg21_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg21_out;
SharedReg28_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg28_out;
SharedReg30_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg30_out;
SharedReg31_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg31_out;
SharedReg34_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg34_out;
SharedReg34_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg34_out;
SharedReg840_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg840_out;
SharedReg551_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg551_out;
SharedReg440_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_13_cast <= SharedReg440_out;
SharedReg441_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_14_cast <= SharedReg441_out;
SharedReg333_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_15_cast <= SharedReg333_out;
SharedReg886_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_16_cast <= SharedReg886_out;
SharedReg551_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_17_cast <= SharedReg551_out;
SharedReg839_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_18_cast <= SharedReg839_out;
SharedReg552_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_19_cast <= SharedReg552_out;
SharedReg882_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_20_cast <= SharedReg882_out;
SharedReg551_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_21_cast <= SharedReg551_out;
SharedReg687_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_22_cast <= SharedReg687_out;
SharedReg551_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_23_cast <= SharedReg551_out;
SharedReg333_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_24_cast <= SharedReg333_out;
SharedReg846_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_25_cast <= SharedReg846_out;
SharedReg551_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_26_cast <= SharedReg551_out;
SharedReg341_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_27_cast <= SharedReg341_out;
SharedReg984_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_28_cast <= SharedReg984_out;
SharedReg556_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_29_cast <= SharedReg556_out;
SharedReg558_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_30_cast <= SharedReg558_out;
SharedReg207_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_31_cast <= SharedReg207_out;
SharedReg447_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_32_cast <= SharedReg447_out;
Delay78No6_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_33_cast <= Delay78No6_out;
SharedReg163_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_34_cast <= SharedReg163_out;
SharedReg853_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_35_cast <= SharedReg853_out;
SharedReg553_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_36_cast <= SharedReg553_out;
Delay44No6_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_37_cast <= Delay44No6_out;
SharedReg844_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_38_cast <= SharedReg844_out;
SharedReg345_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_39_cast <= SharedReg345_out;
SharedReg841_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_40_cast <= SharedReg841_out;
SharedReg1000_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_41_cast <= SharedReg1000_out;
SharedReg188_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_42_cast <= SharedReg188_out;
SharedReg822_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_43_cast <= SharedReg822_out;
SharedReg553_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_44_cast <= SharedReg553_out;
SharedReg842_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_45_cast <= SharedReg842_out;
SharedReg984_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_46_cast <= SharedReg984_out;
SharedReg163_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_47_cast <= SharedReg163_out;
   MUX_Subtract3_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_47_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg25_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg18_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg840_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg551_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg440_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg441_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg333_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg886_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg551_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg839_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg552_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg882_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg19_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg551_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg687_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg551_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg333_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg846_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg551_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg341_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg984_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg556_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg558_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg21_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg207_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg447_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => Delay78No6_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg163_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg853_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg553_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => Delay44No6_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg844_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg345_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg841_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg21_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg1000_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg188_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg822_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg553_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg842_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg984_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg163_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_47_cast,
                 iS_5 => SharedReg28_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg30_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg31_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg34_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg34_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Subtract3_6_impl_1_LUT_out,
                 oMux => MUX_Subtract3_6_impl_1_out);

   Delay1No117_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_6_impl_1_out,
                 Y => Delay1No117_out);

Delay1No118_out_to_Subtract6_2_impl_parent_implementedSystem_port_0_cast <= Delay1No118_out;
Delay1No119_out_to_Subtract6_2_impl_parent_implementedSystem_port_1_cast <= Delay1No119_out;
   Subtract6_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract6_2_impl_out,
                 X => Delay1No118_out_to_Subtract6_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No119_out_to_Subtract6_2_impl_parent_implementedSystem_port_1_cast);

SharedReg237_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg237_out;
SharedReg380_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg380_out;
SharedReg92_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg92_out;
SharedReg380_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg380_out;
SharedReg382_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg382_out;
SharedReg487_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg487_out;
SharedReg599_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg599_out;
SharedReg382_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg382_out;
SharedReg380_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg380_out;
SharedReg747_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg747_out;
SharedReg1_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1_out;
SharedReg3_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg3_out;
SharedReg17_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg17_out;
SharedReg6_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg6_out;
SharedReg11_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg11_out;
SharedReg12_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg12_out;
SharedReg16_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg16_out;
SharedReg380_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg380_out;
SharedReg477_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg477_out;
SharedReg474_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg474_out;
SharedReg71_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg71_out;
SharedReg602_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg602_out;
SharedReg759_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg759_out;
SharedReg377_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg377_out;
SharedReg474_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg474_out;
SharedReg374_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg374_out;
SharedReg8_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg8_out;
SharedReg225_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg225_out;
SharedReg974_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_29_cast <= SharedReg974_out;
SharedReg974_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_30_cast <= SharedReg974_out;
SharedReg236_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_31_cast <= SharedReg236_out;
SharedReg595_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_32_cast <= SharedReg595_out;
SharedReg747_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_33_cast <= SharedReg747_out;
SharedReg82_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_34_cast <= SharedReg82_out;
SharedReg597_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_35_cast <= SharedReg597_out;
SharedReg471_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_36_cast <= SharedReg471_out;
SharedReg239_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_37_cast <= SharedReg239_out;
SharedReg747_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_38_cast <= SharedReg747_out;
SharedReg68_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_39_cast <= SharedReg68_out;
SharedReg933_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_40_cast <= SharedReg933_out;
SharedReg619_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_41_cast <= SharedReg619_out;
SharedReg381_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_42_cast <= SharedReg381_out;
SharedReg603_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_43_cast <= SharedReg603_out;
SharedReg602_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_44_cast <= SharedReg602_out;
SharedReg76_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_45_cast <= SharedReg76_out;
SharedReg605_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_46_cast <= SharedReg605_out;
SharedReg477_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_47_cast <= SharedReg477_out;
SharedReg368_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_48_cast <= SharedReg368_out;
SharedReg617_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_49_cast <= SharedReg617_out;
SharedReg942_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_50_cast <= SharedReg942_out;
SharedReg272_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_51_cast <= SharedReg272_out;
SharedReg79_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_52_cast <= SharedReg79_out;
SharedReg594_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_53_cast <= SharedReg594_out;
SharedReg236_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_54_cast <= SharedReg236_out;
SharedReg103_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_55_cast <= SharedReg103_out;
SharedReg384_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_56_cast <= SharedReg384_out;
SharedReg491_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_57_cast <= SharedReg491_out;
SharedReg490_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_58_cast <= SharedReg490_out;
SharedReg395_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_59_cast <= SharedReg395_out;
SharedReg935_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_60_cast <= SharedReg935_out;
SharedReg766_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_61_cast <= SharedReg766_out;
SharedReg634_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_62_cast <= SharedReg634_out;
SharedReg381_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_63_cast <= SharedReg381_out;
SharedReg908_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_64_cast <= SharedReg908_out;
   MUX_Subtract6_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg237_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg380_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg3_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg17_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg6_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg11_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg12_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg16_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg380_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg477_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg474_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg92_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg71_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg602_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg759_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg377_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg474_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg374_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg8_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg225_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg974_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg974_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg380_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg236_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg595_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg747_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg82_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg597_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg471_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg239_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg747_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg68_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg933_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg382_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg619_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg381_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg603_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg602_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg76_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg605_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg477_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg368_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg617_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg942_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg487_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg272_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg79_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg594_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg236_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg103_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg384_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg491_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg490_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg395_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg935_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg599_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg766_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg634_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg381_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg908_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg382_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg380_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg747_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract6_2_impl_0_out);

   Delay1No118_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract6_2_impl_0_out,
                 Y => Delay1No118_out);

SharedReg107_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg107_out;
SharedReg488_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg488_out;
SharedReg112_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg112_out;
SharedReg766_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg766_out;
SharedReg487_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg487_out;
SharedReg774_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg774_out;
SharedReg906_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg906_out;
SharedReg768_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg768_out;
SharedReg497_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg497_out;
SharedReg750_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg750_out;
SharedReg19_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg19_out;
SharedReg21_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg21_out;
SharedReg35_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg35_out;
SharedReg24_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg24_out;
SharedReg29_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg30_out;
SharedReg34_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg34_out;
SharedReg489_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg489_out;
SharedReg753_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg753_out;
SharedReg753_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg753_out;
SharedReg72_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg72_out;
SharedReg603_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg603_out;
SharedReg762_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg762_out;
Delay43No8_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_24_cast <= Delay43No8_out;
SharedReg747_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg747_out;
SharedReg372_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg372_out;
SharedReg26_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg26_out;
SharedReg62_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg62_out;
SharedReg907_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_29_cast <= SharedReg907_out;
SharedReg595_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_30_cast <= SharedReg595_out;
SharedReg86_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_31_cast <= SharedReg86_out;
SharedReg929_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_32_cast <= SharedReg929_out;
SharedReg757_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_33_cast <= SharedReg757_out;
SharedReg240_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_34_cast <= SharedReg240_out;
Delay76No1_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_35_cast <= Delay76No1_out;
SharedReg752_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_36_cast <= SharedReg752_out;
Delay77No1_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_37_cast <= Delay77No1_out;
SharedReg753_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_38_cast <= SharedReg753_out;
SharedReg235_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_39_cast <= SharedReg235_out;
SharedReg638_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_40_cast <= SharedReg638_out;
SharedReg955_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_41_cast <= SharedReg955_out;
SharedReg487_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_42_cast <= SharedReg487_out;
SharedReg906_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_43_cast <= SharedReg906_out;
SharedReg593_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_44_cast <= SharedReg593_out;
SharedReg235_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_45_cast <= SharedReg235_out;
SharedReg567_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_46_cast <= SharedReg567_out;
SharedReg482_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_47_cast <= SharedReg482_out;
SharedReg476_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_48_cast <= SharedReg476_out;
SharedReg622_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_49_cast <= SharedReg622_out;
SharedReg617_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_50_cast <= SharedReg617_out;
SharedReg88_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_51_cast <= SharedReg88_out;
SharedReg62_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_52_cast <= SharedReg62_out;
SharedReg612_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_53_cast <= SharedReg612_out;
SharedReg84_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_54_cast <= SharedReg84_out;
SharedReg234_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_55_cast <= SharedReg234_out;
SharedReg781_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_56_cast <= SharedReg781_out;
SharedReg772_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_57_cast <= SharedReg772_out;
SharedReg770_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_58_cast <= SharedReg770_out;
SharedReg405_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_59_cast <= SharedReg405_out;
SharedReg621_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_60_cast <= SharedReg621_out;
SharedReg487_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_61_cast <= SharedReg487_out;
SharedReg618_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_62_cast <= SharedReg618_out;
SharedReg487_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_63_cast <= SharedReg487_out;
SharedReg637_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_64_cast <= SharedReg637_out;
   MUX_Subtract6_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg107_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg488_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg19_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg21_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg35_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg24_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg29_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg30_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg34_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg489_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg753_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg753_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg112_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg72_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg603_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg762_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => Delay43No8_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg747_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg372_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg26_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg62_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg907_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg595_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg766_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg86_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg929_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg757_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg240_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => Delay76No1_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg752_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => Delay77No1_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg753_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg235_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg638_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg487_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg955_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg487_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg906_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg593_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg235_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg567_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg482_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg476_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg622_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg617_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg774_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg88_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg62_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg612_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg84_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg234_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg781_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg772_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg770_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg405_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg621_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg906_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg487_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg618_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg487_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg637_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg768_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg497_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg750_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract6_2_impl_1_out);

   Delay1No119_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract6_2_impl_1_out,
                 Y => Delay1No119_out);

Delay1No120_out_to_Subtract6_4_impl_parent_implementedSystem_port_0_cast <= Delay1No120_out;
Delay1No121_out_to_Subtract6_4_impl_parent_implementedSystem_port_1_cast <= Delay1No121_out;
   Subtract6_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract6_4_impl_out,
                 X => Delay1No120_out_to_Subtract6_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No121_out_to_Subtract6_4_impl_parent_implementedSystem_port_1_cast);

SharedReg399_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg399_out;
SharedReg507_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg507_out;
SharedReg506_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg506_out;
SharedReg410_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg410_out;
SharedReg644_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg644_out;
SharedReg784_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg784_out;
SharedReg946_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg946_out;
SharedReg396_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg396_out;
SharedReg933_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg933_out;
SharedReg263_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg263_out;
SharedReg395_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg395_out;
SharedReg118_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg118_out;
SharedReg395_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg395_out;
SharedReg397_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg397_out;
SharedReg503_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg503_out;
SharedReg623_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg623_out;
SharedReg397_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg397_out;
SharedReg802_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg802_out;
SharedReg765_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg765_out;
SharedReg1_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg1_out;
SharedReg3_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg3_out;
SharedReg17_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg17_out;
SharedReg6_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg6_out;
SharedReg11_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg11_out;
SharedReg12_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg12_out;
SharedReg16_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg16_out;
SharedReg395_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg395_out;
SharedReg493_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg493_out;
SharedReg490_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_29_cast <= SharedReg490_out;
SharedReg96_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_30_cast <= SharedReg96_out;
SharedReg627_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_31_cast <= SharedReg627_out;
SharedReg777_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_32_cast <= SharedReg777_out;
SharedReg392_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_33_cast <= SharedReg392_out;
SharedReg490_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_34_cast <= SharedReg490_out;
SharedReg389_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_35_cast <= SharedReg389_out;
SharedReg8_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_36_cast <= SharedReg8_out;
SharedReg251_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_37_cast <= SharedReg251_out;
SharedReg922_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_38_cast <= SharedReg922_out;
SharedReg922_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_39_cast <= SharedReg922_out;
SharedReg633_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_40_cast <= SharedReg633_out;
SharedReg795_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_41_cast <= SharedReg795_out;
SharedReg503_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_42_cast <= SharedReg503_out;
SharedReg109_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_43_cast <= SharedReg109_out;
SharedReg621_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_44_cast <= SharedReg621_out;
SharedReg487_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_45_cast <= SharedReg487_out;
SharedReg265_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_46_cast <= SharedReg265_out;
SharedReg765_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_47_cast <= SharedReg765_out;
SharedReg93_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_48_cast <= SharedReg93_out;
SharedReg642_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_49_cast <= SharedReg642_out;
SharedReg642_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_50_cast <= SharedReg642_out;
SharedReg783_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_51_cast <= SharedReg783_out;
SharedReg628_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_52_cast <= SharedReg628_out;
SharedReg627_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_53_cast <= SharedReg627_out;
SharedReg101_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_54_cast <= SharedReg101_out;
SharedReg861_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_55_cast <= SharedReg861_out;
SharedReg506_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_56_cast <= SharedReg506_out;
SharedReg503_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_57_cast <= SharedReg503_out;
SharedReg285_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_58_cast <= SharedReg285_out;
SharedReg141_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_59_cast <= SharedReg141_out;
SharedReg411_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_60_cast <= SharedReg411_out;
SharedReg114_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_61_cast <= SharedReg114_out;
SharedReg124_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_62_cast <= SharedReg124_out;
SharedReg933_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_63_cast <= SharedReg933_out;
SharedReg651_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_64_cast <= SharedReg651_out;
   MUX_Subtract6_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg399_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg507_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg395_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg118_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg395_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg397_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg503_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg623_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg397_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg802_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg765_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg1_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg506_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg3_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg17_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg6_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg11_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg12_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg16_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg395_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg493_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg490_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg96_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg410_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg627_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg777_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg392_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg490_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg389_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg8_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg251_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg922_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg922_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg633_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg644_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg795_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg503_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg109_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg621_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg487_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg265_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg765_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg93_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg642_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg642_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg784_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg783_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg628_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg627_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg101_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg861_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg506_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg503_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg285_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg141_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg411_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg946_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg114_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg124_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg933_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg651_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg396_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg933_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg263_out_to_MUX_Subtract6_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract6_4_impl_0_out);

   Delay1No120_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract6_4_impl_0_out,
                 Y => Delay1No120_out);

SharedReg799_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg799_out;
SharedReg790_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg790_out;
SharedReg788_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg788_out;
SharedReg420_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg420_out;
SharedReg935_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg935_out;
SharedReg503_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg503_out;
SharedReg641_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg641_out;
SharedReg503_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg503_out;
SharedReg658_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg658_out;
SharedReg132_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg132_out;
SharedReg504_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg504_out;
SharedReg137_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg137_out;
SharedReg784_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg784_out;
SharedReg503_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg503_out;
SharedReg792_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg792_out;
SharedReg931_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg931_out;
SharedReg786_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg786_out;
SharedReg519_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg519_out;
SharedReg768_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg768_out;
SharedReg19_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg19_out;
SharedReg21_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg21_out;
SharedReg35_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg35_out;
SharedReg24_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg24_out;
SharedReg29_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg30_out;
SharedReg34_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg34_out;
SharedReg505_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg505_out;
SharedReg771_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg771_out;
SharedReg771_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_29_cast <= SharedReg771_out;
SharedReg97_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_30_cast <= SharedReg97_out;
SharedReg628_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_31_cast <= SharedReg628_out;
SharedReg780_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_32_cast <= SharedReg780_out;
Delay43No9_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_33_cast <= Delay43No9_out;
SharedReg765_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_34_cast <= SharedReg765_out;
SharedReg387_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_35_cast <= SharedReg387_out;
SharedReg26_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_36_cast <= SharedReg26_out;
SharedReg88_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_37_cast <= SharedReg88_out;
SharedReg932_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_38_cast <= SharedReg932_out;
SharedReg619_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_39_cast <= SharedReg619_out;
SharedReg653_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_40_cast <= SharedReg653_out;
SharedReg798_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_41_cast <= SharedReg798_out;
SharedReg785_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_42_cast <= SharedReg785_out;
SharedReg266_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_43_cast <= SharedReg266_out;
Delay76No2_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_44_cast <= Delay76No2_out;
SharedReg770_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_45_cast <= SharedReg770_out;
Delay77No2_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_46_cast <= Delay77No2_out;
SharedReg771_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_47_cast <= SharedReg771_out;
SharedReg89_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_48_cast <= SharedReg89_out;
SharedReg659_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_49_cast <= SharedReg659_out;
SharedReg880_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_50_cast <= SharedReg880_out;
SharedReg793_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_51_cast <= SharedReg793_out;
SharedReg931_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_52_cast <= SharedReg931_out;
SharedReg617_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_53_cast <= SharedReg617_out;
SharedReg261_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_54_cast <= SharedReg261_out;
Delay78No3_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_55_cast <= Delay78No3_out;
SharedReg503_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_56_cast <= SharedReg503_out;
SharedReg785_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_57_cast <= SharedReg785_out;
SharedReg291_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_58_cast <= SharedReg291_out;
SharedReg330_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_59_cast <= SharedReg330_out;
SharedReg519_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_60_cast <= SharedReg519_out;
SharedReg287_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_61_cast <= SharedReg287_out;
SharedReg260_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_62_cast <= SharedReg260_out;
SharedReg859_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_63_cast <= SharedReg859_out;
SharedReg906_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_64_cast <= SharedReg906_out;
   MUX_Subtract6_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg799_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg790_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg504_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg137_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg784_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg503_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg792_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg931_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg786_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg519_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg768_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg19_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg788_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg21_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg35_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg24_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg29_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg30_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg34_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg505_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg771_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg771_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg97_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg420_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg628_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg780_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => Delay43No9_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg765_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg387_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg26_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg88_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg932_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg619_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg653_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg935_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg798_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg785_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg266_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => Delay76No2_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg770_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => Delay77No2_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg771_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg89_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg659_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg880_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg503_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg793_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg931_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg617_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg261_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => Delay78No3_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg503_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg785_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg291_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg330_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg519_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg641_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg287_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg260_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg859_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg906_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg503_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg658_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg132_out_to_MUX_Subtract6_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract6_4_impl_1_out);

   Delay1No121_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract6_4_impl_1_out,
                 Y => Delay1No121_out);

Delay1No122_out_to_Subtract10_1_impl_parent_implementedSystem_port_0_cast <= Delay1No122_out;
Delay1No123_out_to_Subtract10_1_impl_parent_implementedSystem_port_1_cast <= Delay1No123_out;
   Subtract10_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract10_1_impl_out,
                 X => Delay1No122_out_to_Subtract10_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No123_out_to_Subtract10_1_impl_parent_implementedSystem_port_1_cast);

SharedReg729_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg729_out;
SharedReg1_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1_out;
SharedReg3_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg3_out;
SharedReg17_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg17_out;
SharedReg6_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg6_out;
SharedReg11_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg11_out;
SharedReg12_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg12_out;
SharedReg16_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg16_out;
SharedReg13_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg13_out;
SharedReg461_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg461_out;
SharedReg458_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg458_out;
SharedReg45_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg45_out;
SharedReg576_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg576_out;
SharedReg741_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg741_out;
SharedReg362_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg362_out;
SharedReg458_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg458_out;
SharedReg359_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg359_out;
SharedReg8_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg8_out;
SharedReg55_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg55_out;
SharedReg585_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg585_out;
SharedReg585_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg585_out;
SharedReg210_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg210_out;
SharedReg569_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg569_out;
SharedReg729_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg729_out;
SharedReg230_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg230_out;
SharedReg571_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg571_out;
SharedReg455_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg455_out;
SharedReg213_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg213_out;
SharedReg729_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_29_cast <= SharedReg729_out;
SharedReg214_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_30_cast <= SharedReg214_out;
SharedReg208_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_31_cast <= SharedReg208_out;
SharedReg968_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_32_cast <= SharedReg968_out;
SharedReg220_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_33_cast <= SharedReg220_out;
SharedReg577_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_34_cast <= SharedReg577_out;
SharedReg576_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_35_cast <= SharedReg576_out;
SharedReg50_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_36_cast <= SharedReg50_out;
SharedReg579_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_37_cast <= SharedReg579_out;
SharedReg461_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_38_cast <= SharedReg461_out;
SharedReg353_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_39_cast <= SharedReg353_out;
SharedReg593_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_40_cast <= SharedReg593_out;
SharedReg917_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_41_cast <= SharedReg917_out;
SharedReg910_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_42_cast <= SharedReg910_out;
SharedReg54_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_43_cast <= SharedReg54_out;
SharedReg568_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_44_cast <= SharedReg568_out;
SharedReg210_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_45_cast <= SharedReg210_out;
SharedReg569_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_46_cast <= SharedReg569_out;
SharedReg960_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_47_cast <= SharedReg960_out;
SharedReg462_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_48_cast <= SharedReg462_out;
SharedReg571_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_49_cast <= SharedReg571_out;
SharedReg41_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_50_cast <= SharedReg41_out;
SharedReg366_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_51_cast <= SharedReg366_out;
SharedReg41_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_52_cast <= SharedReg41_out;
SharedReg213_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_53_cast <= SharedReg213_out;
SharedReg573_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_54_cast <= SharedReg573_out;
SharedReg748_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_55_cast <= SharedReg748_out;
SharedReg65_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_56_cast <= SharedReg65_out;
SharedReg365_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_57_cast <= SharedReg365_out;
SharedReg239_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_58_cast <= SharedReg239_out;
SharedReg365_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_59_cast <= SharedReg365_out;
SharedReg367_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_60_cast <= SharedReg367_out;
SharedReg471_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_61_cast <= SharedReg471_out;
SharedReg963_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_62_cast <= SharedReg963_out;
SharedReg367_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_63_cast <= SharedReg367_out;
SharedReg365_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_64_cast <= SharedReg365_out;
   MUX_Subtract10_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg729_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg458_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg45_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg576_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg741_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg362_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg458_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg359_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg8_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg55_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg585_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg3_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg585_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg210_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg569_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg729_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg230_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg571_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg455_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg213_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg729_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg214_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg17_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg208_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg968_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg220_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg577_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg576_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg50_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg579_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg461_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg353_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg593_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg6_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg917_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg910_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg54_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg568_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg210_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg569_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg960_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg462_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg571_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg41_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg11_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg366_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg41_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg213_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg573_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg748_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg65_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg365_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg239_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg365_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg367_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg12_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg471_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg963_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg367_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg365_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg16_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg13_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg461_out_to_MUX_Subtract10_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract10_1_impl_0_out);

   Delay1No122_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract10_1_impl_0_out,
                 Y => Delay1No122_out);

SharedReg732_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg732_out;
SharedReg19_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg19_out;
SharedReg21_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg21_out;
SharedReg35_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg35_out;
SharedReg24_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg24_out;
SharedReg29_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg30_out;
SharedReg34_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg34_out;
SharedReg31_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg31_out;
SharedReg735_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg735_out;
SharedReg735_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg735_out;
SharedReg46_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg46_out;
SharedReg577_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg577_out;
SharedReg744_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg744_out;
Delay43No7_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_15_cast <= Delay43No7_out;
SharedReg729_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg729_out;
SharedReg357_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg357_out;
SharedReg26_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg26_out;
SharedReg36_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg36_out;
SharedReg958_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg958_out;
SharedReg569_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg569_out;
SharedReg60_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg60_out;
SharedReg981_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg981_out;
SharedReg739_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg739_out;
SharedReg214_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg214_out;
Delay76No_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_26_cast <= Delay76No_out;
SharedReg734_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg734_out;
Delay77No_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_28_cast <= Delay77No_out;
SharedReg735_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_29_cast <= SharedReg735_out;
SharedReg209_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_30_cast <= SharedReg209_out;
SharedReg214_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_31_cast <= SharedReg214_out;
SharedReg567_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_32_cast <= SharedReg567_out;
SharedReg36_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_33_cast <= SharedReg36_out;
SharedReg957_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_34_cast <= SharedReg957_out;
SharedReg567_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_35_cast <= SharedReg567_out;
SharedReg209_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_36_cast <= SharedReg209_out;
SharedReg567_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_37_cast <= SharedReg567_out;
SharedReg466_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_38_cast <= SharedReg466_out;
SharedReg460_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_39_cast <= SharedReg460_out;
SharedReg598_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_40_cast <= SharedReg598_out;
SharedReg593_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_41_cast <= SharedReg593_out;
SharedReg597_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_42_cast <= SharedReg597_out;
SharedReg36_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_43_cast <= SharedReg36_out;
SharedReg588_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_44_cast <= SharedReg588_out;
SharedReg58_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_45_cast <= SharedReg58_out;
SharedReg588_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_46_cast <= SharedReg588_out;
SharedReg589_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_47_cast <= SharedReg589_out;
SharedReg729_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_48_cast <= SharedReg729_out;
SharedReg980_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_49_cast <= SharedReg980_out;
SharedReg231_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_50_cast <= SharedReg231_out;
SharedReg471_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_51_cast <= SharedReg471_out;
SharedReg208_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_52_cast <= SharedReg208_out;
SharedReg208_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_53_cast <= SharedReg208_out;
SharedReg958_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_54_cast <= SharedReg958_out;
SharedReg471_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_55_cast <= SharedReg471_out;
SharedReg254_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_56_cast <= SharedReg254_out;
SharedReg472_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_57_cast <= SharedReg472_out;
SharedReg85_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_58_cast <= SharedReg85_out;
SharedReg748_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_59_cast <= SharedReg748_out;
SharedReg471_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_60_cast <= SharedReg471_out;
SharedReg756_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_61_cast <= SharedReg756_out;
SharedReg957_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_62_cast <= SharedReg957_out;
SharedReg750_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_63_cast <= SharedReg750_out;
SharedReg481_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_64_cast <= SharedReg481_out;
   MUX_Subtract10_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_64_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg732_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg19_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg735_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg46_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg577_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg744_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => Delay43No7_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg729_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg357_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg26_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg36_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg958_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg21_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg569_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg60_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg981_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg739_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg214_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => Delay76No_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg734_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => Delay77No_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg735_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg209_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg35_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg214_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg567_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg36_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg957_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg567_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg209_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg567_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg466_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg460_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg598_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg24_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg593_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg597_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg36_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg588_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg58_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg588_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg589_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg729_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg980_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg231_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg29_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg471_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg208_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg208_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg958_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg471_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg254_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg472_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg85_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg748_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_59_cast,
                 iS_59 => SharedReg471_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_60_cast,
                 iS_6 => SharedReg30_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_60 => SharedReg756_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_61_cast,
                 iS_61 => SharedReg957_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_62_cast,
                 iS_62 => SharedReg750_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_63_cast,
                 iS_63 => SharedReg481_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_64_cast,
                 iS_7 => SharedReg34_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg31_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg735_out_to_MUX_Subtract10_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount641_out,
                 oMux => MUX_Subtract10_1_impl_1_out);

   Delay1No123_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract10_1_impl_1_out,
                 Y => Delay1No123_out);

Delay1No124_out_to_Subtract12_6_impl_parent_implementedSystem_port_0_cast <= Delay1No124_out;
Delay1No125_out_to_Subtract12_6_impl_parent_implementedSystem_port_1_cast <= Delay1No125_out;
   Subtract12_6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract12_6_impl_out,
                 X => Delay1No124_out_to_Subtract12_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No125_out_to_Subtract12_6_impl_parent_implementedSystem_port_1_cast);

SharedReg1_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1_out;
SharedReg11_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg11_out;
SharedReg12_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg12_out;
SharedReg717_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg717_out;
SharedReg891_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg891_out;
SharedReg203_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg203_out;
SharedReg894_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg894_out;
SharedReg177_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg177_out;
SharedReg191_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg191_out;
SharedReg440_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg440_out;
SharedReg442_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg442_out;
SharedReg445_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg445_out;
SharedReg337_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_13_cast <= SharedReg337_out;
SharedReg180_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_14_cast <= SharedReg180_out;
SharedReg699_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_15_cast <= SharedReg699_out;
SharedReg888_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_16_cast <= SharedReg888_out;
SharedReg843_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_17_cast <= SharedReg843_out;
SharedReg558_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_18_cast <= SharedReg558_out;
SharedReg452_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_19_cast <= SharedReg452_out;
SharedReg886_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_20_cast <= SharedReg886_out;
SharedReg168_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_21_cast <= SharedReg168_out;
SharedReg449_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_22_cast <= SharedReg449_out;
SharedReg557_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_23_cast <= SharedReg557_out;
SharedReg554_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_24_cast <= SharedReg554_out;
SharedReg883_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_25_cast <= SharedReg883_out;
SharedReg837_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_26_cast <= SharedReg837_out;
SharedReg884_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_27_cast <= SharedReg884_out;
SharedReg443_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_28_cast <= SharedReg443_out;
SharedReg986_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_29_cast <= SharedReg986_out;
SharedReg837_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_30_cast <= SharedReg837_out;
SharedReg557_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_31_cast <= SharedReg557_out;
SharedReg342_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_32_cast <= SharedReg342_out;
SharedReg554_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_33_cast <= SharedReg554_out;
SharedReg837_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_34_cast <= SharedReg837_out;
   MUX_Subtract12_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_34_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg11_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg442_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg445_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg337_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg180_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg699_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg888_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg843_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg558_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg452_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg886_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg12_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg168_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg449_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg557_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg554_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg883_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg837_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg884_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg443_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg986_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg837_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg717_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg557_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg342_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg554_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg837_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_34_cast,
                 iS_4 => SharedReg891_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg203_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg894_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg177_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg191_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg440_out_to_MUX_Subtract12_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Subtract12_6_impl_0_LUT_out,
                 oMux => MUX_Subtract12_6_impl_0_out);

   Delay1No124_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_6_impl_0_out,
                 Y => Delay1No124_out);

SharedReg19_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg19_out;
SharedReg29_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg30_out;
SharedReg186_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg186_out;
SharedReg186_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg186_out;
SharedReg685_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg685_out;
SharedReg561_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg551_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg551_out;
SharedReg332_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg332_out;
SharedReg564_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg564_out;
SharedReg310_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg310_out;
SharedReg708_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg708_out;
SharedReg169_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_13_cast <= SharedReg169_out;
SharedReg882_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_14_cast <= SharedReg882_out;
SharedReg841_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_15_cast <= SharedReg841_out;
SharedReg332_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_16_cast <= SharedReg332_out;
SharedReg837_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_17_cast <= SharedReg837_out;
Delay43No13_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_18_cast <= Delay43No13_out;
SharedReg447_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_19_cast <= SharedReg447_out;
Delay76No6_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_20_cast <= Delay76No6_out;
Delay77No6_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_21_cast <= Delay77No6_out;
SharedReg843_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_22_cast <= SharedReg843_out;
SharedReg843_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_23_cast <= SharedReg843_out;
SharedReg900_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_24_cast <= SharedReg900_out;
SharedReg843_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_25_cast <= SharedReg843_out;
SharedReg983_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_26_cast <= SharedReg983_out;
SharedReg900_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_27_cast <= SharedReg900_out;
SharedReg556_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_28_cast <= SharedReg556_out;
SharedReg840_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_29_cast <= SharedReg840_out;
SharedReg902_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_30_cast <= SharedReg902_out;
SharedReg707_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_31_cast <= SharedReg707_out;
SharedReg562_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_32_cast <= SharedReg562_out;
SharedReg847_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_33_cast <= SharedReg847_out;
SharedReg837_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_34_cast <= SharedReg837_out;
   MUX_Subtract12_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_34_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg19_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg29_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg310_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg708_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg169_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg882_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg841_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg332_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg837_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => Delay43No13_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg447_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => Delay76No6_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg30_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => Delay77No6_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg843_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg843_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg900_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg843_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg983_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg900_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg556_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg840_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg902_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg186_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg707_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg562_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg847_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg837_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_34_cast,
                 iS_4 => SharedReg186_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg685_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg551_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg332_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg564_out_to_MUX_Subtract12_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Subtract12_6_impl_1_LUT_out,
                 oMux => MUX_Subtract12_6_impl_1_out);

   Delay1No125_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_6_impl_1_out,
                 Y => Delay1No125_out);
   Constant2_0_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant2_0_impl_out);
   Constant11_0_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant11_0_impl_out);
   Constant4_0_impl_instance: Constant_float_8_23_cosnpi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant4_0_impl_out);
   Constant13_0_impl_instance: Constant_float_8_23_sinnpi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant13_0_impl_out);
   Constant5_0_impl_instance: Constant_float_8_23_cosn3_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant5_0_impl_out);
   Constant14_0_impl_instance: Constant_float_8_23_sinn3_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant14_0_impl_out);
   Constant6_0_impl_instance: Constant_float_8_23_cosnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant6_0_impl_out);
   Constant15_0_impl_instance: Constant_float_8_23_sinnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant15_0_impl_out);
   Constant7_0_impl_instance: Constant_float_8_23_cosn5_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant7_0_impl_out);
   Constant16_0_impl_instance: Constant_float_8_23_sinn5_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant16_0_impl_out);
   Constant8_0_impl_instance: Constant_float_8_23_cosn3_mult_pi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant8_0_impl_out);
   Constant17_0_impl_instance: Constant_float_8_23_sinn3_mult_pi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant17_0_impl_out);
   Constant9_0_impl_instance: Constant_float_8_23_cosn7_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant9_0_impl_out);
   Constant18_0_impl_instance: Constant_float_8_23_sinn7_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant18_0_impl_out);
   Constant_0_impl_instance: Constant_float_8_23_cosnpi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant_0_impl_out);
   Constant1_0_impl_instance: Constant_float_8_23_sinnpi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant1_0_impl_out);

   Delay43No_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg364_out,
                 Y => Delay43No_out);

   Delay43No1_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg379_out,
                 Y => Delay43No1_out);

   Delay43No2_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg394_out,
                 Y => Delay43No2_out);

   Delay43No3_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg409_out,
                 Y => Delay43No3_out);

   Delay43No4_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg424_out,
                 Y => Delay43No4_out);

   Delay43No5_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg439_out,
                 Y => Delay43No5_out);

   Delay43No6_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg454_out,
                 Y => Delay43No6_out);

   Delay43No7_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg470_out,
                 Y => Delay43No7_out);

   Delay43No8_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg486_out,
                 Y => Delay43No8_out);

   Delay43No9_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg502_out,
                 Y => Delay43No9_out);

   Delay43No10_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg518_out,
                 Y => Delay43No10_out);

   Delay43No11_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg534_out,
                 Y => Delay43No11_out);

   Delay43No12_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg550_out,
                 Y => Delay43No12_out);

   Delay43No13_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg566_out,
                 Y => Delay43No13_out);

   Delay76No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg592_out,
                 Y => Delay76No_out);

   Delay76No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg616_out,
                 Y => Delay76No1_out);

   Delay76No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg639_out,
                 Y => Delay76No2_out);

   Delay76No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg660_out,
                 Y => Delay76No3_out);

   Delay76No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg684_out,
                 Y => Delay76No4_out);

   Delay76No6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg905_out,
                 Y => Delay76No6_out);

   Delay77No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg233_out,
                 Y => Delay77No_out);

   Delay77No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg259_out,
                 Y => Delay77No1_out);

   Delay77No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg284_out,
                 Y => Delay77No2_out);

   Delay77No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg309_out,
                 Y => Delay77No3_out);

   Delay77No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg331_out,
                 Y => Delay77No4_out);

   Delay77No5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg185_out,
                 Y => Delay77No5_out);

   Delay77No6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg349_out,
                 Y => Delay77No6_out);

   Delay78No_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg982_out,
                 Y => Delay78No_out);

   Delay78No1_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg930_out,
                 Y => Delay78No1_out);

   Delay78No2_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg956_out,
                 Y => Delay78No2_out);

   Delay78No3_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg881_out,
                 Y => Delay78No3_out);

   Delay78No4_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg706_out,
                 Y => Delay78No4_out);

   Delay78No5_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg728_out,
                 Y => Delay78No5_out);

   Delay78No6_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1002_out,
                 Y => Delay78No6_out);

   Delay44No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg746_out,
                 Y => Delay44No_out);

   Delay44No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg764_out,
                 Y => Delay44No1_out);

   Delay44No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg782_out,
                 Y => Delay44No2_out);

   Delay44No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg800_out,
                 Y => Delay44No3_out);

   Delay44No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg818_out,
                 Y => Delay44No4_out);

   Delay44No5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg836_out,
                 Y => Delay44No5_out);

   Delay44No6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg854_out,
                 Y => Delay44No6_out);

   MUX_y0_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y0_re_0_0_LUT_out);

   MUX_y0_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y0_im_0_0_LUT_out);

   MUX_y1_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y1_re_0_0_LUT_out);

   MUX_y1_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y1_im_0_0_LUT_out);

   MUX_y2_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y2_re_0_0_LUT_out);

   MUX_y2_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y2_im_0_0_LUT_out);

   MUX_y3_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y3_re_0_0_LUT_out);

   MUX_y3_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y3_im_0_0_LUT_out);

   MUX_y4_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y4_re_0_0_LUT_out);

   MUX_y4_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y4_im_0_0_LUT_out);

   MUX_y5_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y5_re_0_0_LUT_out);

   MUX_y5_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y5_im_0_0_LUT_out);

   MUX_y6_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y6_re_0_0_LUT_out);

   MUX_y6_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y6_im_0_0_LUT_out);

   MUX_y7_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y7_re_0_0_LUT_out);

   MUX_y7_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y7_im_0_0_LUT_out);

   MUX_y8_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y8_re_0_0_LUT_out);

   MUX_y8_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y8_im_0_0_LUT_out);

   MUX_y9_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y9_re_0_0_LUT_out);

   MUX_y9_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y9_im_0_0_LUT_out);

   MUX_y10_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y10_re_0_0_LUT_out);

   MUX_y10_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y10_im_0_0_LUT_out);

   MUX_y11_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y11_re_0_0_LUT_out);

   MUX_y11_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y11_im_0_0_LUT_out);

   MUX_y12_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y12_re_0_0_LUT_out);

   MUX_y12_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y12_im_0_0_LUT_out);

   MUX_y13_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y13_re_0_0_LUT_out);

   MUX_y13_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y13_im_0_0_LUT_out);

   MUX_y14_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y14_re_0_0_LUT_out);

   MUX_y14_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y14_im_0_0_LUT_out);

   MUX_y15_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y15_re_0_0_LUT_out);

   MUX_y15_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_y15_im_0_0_LUT_out);

   MUX_Add2_5_impl_0_LUT_instance: GenericLut_LUTData_MUX_Add2_5_impl_0_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_Add2_5_impl_0_LUT_out);

   MUX_Add2_5_impl_1_LUT_instance: GenericLut_LUTData_MUX_Add2_5_impl_1_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_Add2_5_impl_1_LUT_out);

   MUX_Add2_6_impl_0_LUT_instance: GenericLut_LUTData_MUX_Add2_6_impl_0_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_Add2_6_impl_0_LUT_out);

   MUX_Add2_6_impl_1_LUT_instance: GenericLut_LUTData_MUX_Add2_6_impl_1_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_Add2_6_impl_1_LUT_out);

   MUX_Add11_6_impl_0_LUT_instance: GenericLut_LUTData_MUX_Add11_6_impl_0_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_Add11_6_impl_0_LUT_out);

   MUX_Add11_6_impl_1_LUT_instance: GenericLut_LUTData_MUX_Add11_6_impl_1_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_Add11_6_impl_1_LUT_out);

   MUX_Subtract2_6_impl_0_LUT_instance: GenericLut_LUTData_MUX_Subtract2_6_impl_0_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_Subtract2_6_impl_0_LUT_out);

   MUX_Subtract2_6_impl_1_LUT_instance: GenericLut_LUTData_MUX_Subtract2_6_impl_1_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_Subtract2_6_impl_1_LUT_out);

   MUX_Subtract3_6_impl_0_LUT_instance: GenericLut_LUTData_MUX_Subtract3_6_impl_0_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_Subtract3_6_impl_0_LUT_out);

   MUX_Subtract3_6_impl_1_LUT_instance: GenericLut_LUTData_MUX_Subtract3_6_impl_1_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_Subtract3_6_impl_1_LUT_out);

   MUX_Subtract12_6_impl_0_LUT_instance: GenericLut_LUTData_MUX_Subtract12_6_impl_0_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_Subtract12_6_impl_0_LUT_out);

   MUX_Subtract12_6_impl_1_LUT_instance: GenericLut_LUTData_MUX_Subtract12_6_impl_1_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount641_out,
                 Output => MUX_Subtract12_6_impl_1_LUT_out);

   SharedReg_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x0_re_0_out,
                 Y => SharedReg_out);

   SharedReg1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x0_im_0_out,
                 Y => SharedReg1_out);

   SharedReg2_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x1_re_0_out,
                 Y => SharedReg2_out);

   SharedReg3_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x1_im_0_out,
                 Y => SharedReg3_out);

   SharedReg4_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x2_re_0_out,
                 Y => SharedReg4_out);

   SharedReg5_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x2_im_0_out,
                 Y => SharedReg5_out);

   SharedReg6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg5_out,
                 Y => SharedReg6_out);

   SharedReg7_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x3_re_0_out,
                 Y => SharedReg7_out);

   SharedReg8_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x3_im_0_out,
                 Y => SharedReg8_out);

   SharedReg9_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x4_re_0_out,
                 Y => SharedReg9_out);

   SharedReg10_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x4_im_0_out,
                 Y => SharedReg10_out);

   SharedReg11_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x5_re_0_out,
                 Y => SharedReg11_out);

   SharedReg12_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x5_im_0_out,
                 Y => SharedReg12_out);

   SharedReg13_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x6_re_0_out,
                 Y => SharedReg13_out);

   SharedReg14_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x6_im_0_out,
                 Y => SharedReg14_out);

   SharedReg15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg14_out,
                 Y => SharedReg15_out);

   SharedReg16_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x7_re_0_out,
                 Y => SharedReg16_out);

   SharedReg17_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x7_im_0_out,
                 Y => SharedReg17_out);

   SharedReg18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x8_re_0_out,
                 Y => SharedReg18_out);

   SharedReg19_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x8_im_0_out,
                 Y => SharedReg19_out);

   SharedReg20_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x9_re_0_out,
                 Y => SharedReg20_out);

   SharedReg21_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x9_im_0_out,
                 Y => SharedReg21_out);

   SharedReg22_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x10_re_0_out,
                 Y => SharedReg22_out);

   SharedReg23_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x10_im_0_out,
                 Y => SharedReg23_out);

   SharedReg24_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg23_out,
                 Y => SharedReg24_out);

   SharedReg25_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x11_re_0_out,
                 Y => SharedReg25_out);

   SharedReg26_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x11_im_0_out,
                 Y => SharedReg26_out);

   SharedReg27_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x12_re_0_out,
                 Y => SharedReg27_out);

   SharedReg28_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x12_im_0_out,
                 Y => SharedReg28_out);

   SharedReg29_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x13_re_0_out,
                 Y => SharedReg29_out);

   SharedReg30_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x13_im_0_out,
                 Y => SharedReg30_out);

   SharedReg31_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x14_re_0_out,
                 Y => SharedReg31_out);

   SharedReg32_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x14_im_0_out,
                 Y => SharedReg32_out);

   SharedReg33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg32_out,
                 Y => SharedReg33_out);

   SharedReg34_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x15_re_0_out,
                 Y => SharedReg34_out);

   SharedReg35_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x15_im_0_out,
                 Y => SharedReg35_out);

   SharedReg36_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_0_impl_out,
                 Y => SharedReg36_out);

   SharedReg37_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg36_out,
                 Y => SharedReg37_out);

   SharedReg38_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg37_out,
                 Y => SharedReg38_out);

   SharedReg39_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg38_out,
                 Y => SharedReg39_out);

   SharedReg40_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg39_out,
                 Y => SharedReg40_out);

   SharedReg41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg40_out,
                 Y => SharedReg41_out);

   SharedReg42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg41_out,
                 Y => SharedReg42_out);

   SharedReg43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg42_out,
                 Y => SharedReg43_out);

   SharedReg44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg43_out,
                 Y => SharedReg44_out);

   SharedReg45_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg44_out,
                 Y => SharedReg45_out);

   SharedReg46_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg45_out,
                 Y => SharedReg46_out);

   SharedReg47_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg46_out,
                 Y => SharedReg47_out);

   SharedReg48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg47_out,
                 Y => SharedReg48_out);

   SharedReg49_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg48_out,
                 Y => SharedReg49_out);

   SharedReg50_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg49_out,
                 Y => SharedReg50_out);

   SharedReg51_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg50_out,
                 Y => SharedReg51_out);

   SharedReg52_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg51_out,
                 Y => SharedReg52_out);

   SharedReg53_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg52_out,
                 Y => SharedReg53_out);

   SharedReg54_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg53_out,
                 Y => SharedReg54_out);

   SharedReg55_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg54_out,
                 Y => SharedReg55_out);

   SharedReg56_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg55_out,
                 Y => SharedReg56_out);

   SharedReg57_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg56_out,
                 Y => SharedReg57_out);

   SharedReg58_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg57_out,
                 Y => SharedReg58_out);

   SharedReg59_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg58_out,
                 Y => SharedReg59_out);

   SharedReg60_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg59_out,
                 Y => SharedReg60_out);

   SharedReg61_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg60_out,
                 Y => SharedReg61_out);

   SharedReg62_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_1_impl_out,
                 Y => SharedReg62_out);

   SharedReg63_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg62_out,
                 Y => SharedReg63_out);

   SharedReg64_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg63_out,
                 Y => SharedReg64_out);

   SharedReg65_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg64_out,
                 Y => SharedReg65_out);

   SharedReg66_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg65_out,
                 Y => SharedReg66_out);

   SharedReg67_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg66_out,
                 Y => SharedReg67_out);

   SharedReg68_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg67_out,
                 Y => SharedReg68_out);

   SharedReg69_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg68_out,
                 Y => SharedReg69_out);

   SharedReg70_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg69_out,
                 Y => SharedReg70_out);

   SharedReg71_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg70_out,
                 Y => SharedReg71_out);

   SharedReg72_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg71_out,
                 Y => SharedReg72_out);

   SharedReg73_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg72_out,
                 Y => SharedReg73_out);

   SharedReg74_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg73_out,
                 Y => SharedReg74_out);

   SharedReg75_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg74_out,
                 Y => SharedReg75_out);

   SharedReg76_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg75_out,
                 Y => SharedReg76_out);

   SharedReg77_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg76_out,
                 Y => SharedReg77_out);

   SharedReg78_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg77_out,
                 Y => SharedReg78_out);

   SharedReg79_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg78_out,
                 Y => SharedReg79_out);

   SharedReg80_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg79_out,
                 Y => SharedReg80_out);

   SharedReg81_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg80_out,
                 Y => SharedReg81_out);

   SharedReg82_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg81_out,
                 Y => SharedReg82_out);

   SharedReg83_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg82_out,
                 Y => SharedReg83_out);

   SharedReg84_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg83_out,
                 Y => SharedReg84_out);

   SharedReg85_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg84_out,
                 Y => SharedReg85_out);

   SharedReg86_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg85_out,
                 Y => SharedReg86_out);

   SharedReg87_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg86_out,
                 Y => SharedReg87_out);

   SharedReg88_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_2_impl_out,
                 Y => SharedReg88_out);

   SharedReg89_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg88_out,
                 Y => SharedReg89_out);

   SharedReg90_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg89_out,
                 Y => SharedReg90_out);

   SharedReg91_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg90_out,
                 Y => SharedReg91_out);

   SharedReg92_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg91_out,
                 Y => SharedReg92_out);

   SharedReg93_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg92_out,
                 Y => SharedReg93_out);

   SharedReg94_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg93_out,
                 Y => SharedReg94_out);

   SharedReg95_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg94_out,
                 Y => SharedReg95_out);

   SharedReg96_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg95_out,
                 Y => SharedReg96_out);

   SharedReg97_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg96_out,
                 Y => SharedReg97_out);

   SharedReg98_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg97_out,
                 Y => SharedReg98_out);

   SharedReg99_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg98_out,
                 Y => SharedReg99_out);

   SharedReg100_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg99_out,
                 Y => SharedReg100_out);

   SharedReg101_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg100_out,
                 Y => SharedReg101_out);

   SharedReg102_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg101_out,
                 Y => SharedReg102_out);

   SharedReg103_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg102_out,
                 Y => SharedReg103_out);

   SharedReg104_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg103_out,
                 Y => SharedReg104_out);

   SharedReg105_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg104_out,
                 Y => SharedReg105_out);

   SharedReg106_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg105_out,
                 Y => SharedReg106_out);

   SharedReg107_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg106_out,
                 Y => SharedReg107_out);

   SharedReg108_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg107_out,
                 Y => SharedReg108_out);

   SharedReg109_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg108_out,
                 Y => SharedReg109_out);

   SharedReg110_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg109_out,
                 Y => SharedReg110_out);

   SharedReg111_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg110_out,
                 Y => SharedReg111_out);

   SharedReg112_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg111_out,
                 Y => SharedReg112_out);

   SharedReg113_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg112_out,
                 Y => SharedReg113_out);

   SharedReg114_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_3_impl_out,
                 Y => SharedReg114_out);

   SharedReg115_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg114_out,
                 Y => SharedReg115_out);

   SharedReg116_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg115_out,
                 Y => SharedReg116_out);

   SharedReg117_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg116_out,
                 Y => SharedReg117_out);

   SharedReg118_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg117_out,
                 Y => SharedReg118_out);

   SharedReg119_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg118_out,
                 Y => SharedReg119_out);

   SharedReg120_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg119_out,
                 Y => SharedReg120_out);

   SharedReg121_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg120_out,
                 Y => SharedReg121_out);

   SharedReg122_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg121_out,
                 Y => SharedReg122_out);

   SharedReg123_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg122_out,
                 Y => SharedReg123_out);

   SharedReg124_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg123_out,
                 Y => SharedReg124_out);

   SharedReg125_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg124_out,
                 Y => SharedReg125_out);

   SharedReg126_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg125_out,
                 Y => SharedReg126_out);

   SharedReg127_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg126_out,
                 Y => SharedReg127_out);

   SharedReg128_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg127_out,
                 Y => SharedReg128_out);

   SharedReg129_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg128_out,
                 Y => SharedReg129_out);

   SharedReg130_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg129_out,
                 Y => SharedReg130_out);

   SharedReg131_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg130_out,
                 Y => SharedReg131_out);

   SharedReg132_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg131_out,
                 Y => SharedReg132_out);

   SharedReg133_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg132_out,
                 Y => SharedReg133_out);

   SharedReg134_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg133_out,
                 Y => SharedReg134_out);

   SharedReg135_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg134_out,
                 Y => SharedReg135_out);

   SharedReg136_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg135_out,
                 Y => SharedReg136_out);

   SharedReg137_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg136_out,
                 Y => SharedReg137_out);

   SharedReg138_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg137_out,
                 Y => SharedReg138_out);

   SharedReg139_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_4_impl_out,
                 Y => SharedReg139_out);

   SharedReg140_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg139_out,
                 Y => SharedReg140_out);

   SharedReg141_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg140_out,
                 Y => SharedReg141_out);

   SharedReg142_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg141_out,
                 Y => SharedReg142_out);

   SharedReg143_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg142_out,
                 Y => SharedReg143_out);

   SharedReg144_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg143_out,
                 Y => SharedReg144_out);

   SharedReg145_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg144_out,
                 Y => SharedReg145_out);

   SharedReg146_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg145_out,
                 Y => SharedReg146_out);

   SharedReg147_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg146_out,
                 Y => SharedReg147_out);

   SharedReg148_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg147_out,
                 Y => SharedReg148_out);

   SharedReg149_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg148_out,
                 Y => SharedReg149_out);

   SharedReg150_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg149_out,
                 Y => SharedReg150_out);

   SharedReg151_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg150_out,
                 Y => SharedReg151_out);

   SharedReg152_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg151_out,
                 Y => SharedReg152_out);

   SharedReg153_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg152_out,
                 Y => SharedReg153_out);

   SharedReg154_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg153_out,
                 Y => SharedReg154_out);

   SharedReg155_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg154_out,
                 Y => SharedReg155_out);

   SharedReg156_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg155_out,
                 Y => SharedReg156_out);

   SharedReg157_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg156_out,
                 Y => SharedReg157_out);

   SharedReg158_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg157_out,
                 Y => SharedReg158_out);

   SharedReg159_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg158_out,
                 Y => SharedReg159_out);

   SharedReg160_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg159_out,
                 Y => SharedReg160_out);

   SharedReg161_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg160_out,
                 Y => SharedReg161_out);

   SharedReg162_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg161_out,
                 Y => SharedReg162_out);

   SharedReg163_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_5_impl_out,
                 Y => SharedReg163_out);

   SharedReg164_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg163_out,
                 Y => SharedReg164_out);

   SharedReg165_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg164_out,
                 Y => SharedReg165_out);

   SharedReg166_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg165_out,
                 Y => SharedReg166_out);

   SharedReg167_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg166_out,
                 Y => SharedReg167_out);

   SharedReg168_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg167_out,
                 Y => SharedReg168_out);

   SharedReg169_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg168_out,
                 Y => SharedReg169_out);

   SharedReg170_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg169_out,
                 Y => SharedReg170_out);

   SharedReg171_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg170_out,
                 Y => SharedReg171_out);

   SharedReg172_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg171_out,
                 Y => SharedReg172_out);

   SharedReg173_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg172_out,
                 Y => SharedReg173_out);

   SharedReg174_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg173_out,
                 Y => SharedReg174_out);

   SharedReg175_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg174_out,
                 Y => SharedReg175_out);

   SharedReg176_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg175_out,
                 Y => SharedReg176_out);

   SharedReg177_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg176_out,
                 Y => SharedReg177_out);

   SharedReg178_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg177_out,
                 Y => SharedReg178_out);

   SharedReg179_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg178_out,
                 Y => SharedReg179_out);

   SharedReg180_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg179_out,
                 Y => SharedReg180_out);

   SharedReg181_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg180_out,
                 Y => SharedReg181_out);

   SharedReg182_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg181_out,
                 Y => SharedReg182_out);

   SharedReg183_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg182_out,
                 Y => SharedReg183_out);

   SharedReg184_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg183_out,
                 Y => SharedReg184_out);

   SharedReg185_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg184_out,
                 Y => SharedReg185_out);

   SharedReg186_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_6_impl_out,
                 Y => SharedReg186_out);

   SharedReg187_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg186_out,
                 Y => SharedReg187_out);

   SharedReg188_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg187_out,
                 Y => SharedReg188_out);

   SharedReg189_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg188_out,
                 Y => SharedReg189_out);

   SharedReg190_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg189_out,
                 Y => SharedReg190_out);

   SharedReg191_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg190_out,
                 Y => SharedReg191_out);

   SharedReg192_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg191_out,
                 Y => SharedReg192_out);

   SharedReg193_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg192_out,
                 Y => SharedReg193_out);

   SharedReg194_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg193_out,
                 Y => SharedReg194_out);

   SharedReg195_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg194_out,
                 Y => SharedReg195_out);

   SharedReg196_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg195_out,
                 Y => SharedReg196_out);

   SharedReg197_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg196_out,
                 Y => SharedReg197_out);

   SharedReg198_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg197_out,
                 Y => SharedReg198_out);

   SharedReg199_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg198_out,
                 Y => SharedReg199_out);

   SharedReg200_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg199_out,
                 Y => SharedReg200_out);

   SharedReg201_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg200_out,
                 Y => SharedReg201_out);

   SharedReg202_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg201_out,
                 Y => SharedReg202_out);

   SharedReg203_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg202_out,
                 Y => SharedReg203_out);

   SharedReg204_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg203_out,
                 Y => SharedReg204_out);

   SharedReg205_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg204_out,
                 Y => SharedReg205_out);

   SharedReg206_instance: Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=30 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg205_out,
                 Y => SharedReg206_out);

   SharedReg207_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg206_out,
                 Y => SharedReg207_out);

   SharedReg208_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_0_impl_out,
                 Y => SharedReg208_out);

   SharedReg209_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg208_out,
                 Y => SharedReg209_out);

   SharedReg210_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg209_out,
                 Y => SharedReg210_out);

   SharedReg211_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg210_out,
                 Y => SharedReg211_out);

   SharedReg212_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg211_out,
                 Y => SharedReg212_out);

   SharedReg213_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg212_out,
                 Y => SharedReg213_out);

   SharedReg214_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg213_out,
                 Y => SharedReg214_out);

   SharedReg215_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg214_out,
                 Y => SharedReg215_out);

   SharedReg216_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg215_out,
                 Y => SharedReg216_out);

   SharedReg217_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg216_out,
                 Y => SharedReg217_out);

   SharedReg218_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg217_out,
                 Y => SharedReg218_out);

   SharedReg219_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg218_out,
                 Y => SharedReg219_out);

   SharedReg220_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg219_out,
                 Y => SharedReg220_out);

   SharedReg221_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg220_out,
                 Y => SharedReg221_out);

   SharedReg222_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg221_out,
                 Y => SharedReg222_out);

   SharedReg223_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg222_out,
                 Y => SharedReg223_out);

   SharedReg224_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg223_out,
                 Y => SharedReg224_out);

   SharedReg225_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg224_out,
                 Y => SharedReg225_out);

   SharedReg226_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg225_out,
                 Y => SharedReg226_out);

   SharedReg227_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg226_out,
                 Y => SharedReg227_out);

   SharedReg228_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg227_out,
                 Y => SharedReg228_out);

   SharedReg229_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg228_out,
                 Y => SharedReg229_out);

   SharedReg230_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg229_out,
                 Y => SharedReg230_out);

   SharedReg231_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg230_out,
                 Y => SharedReg231_out);

   SharedReg232_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg231_out,
                 Y => SharedReg232_out);

   SharedReg233_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg232_out,
                 Y => SharedReg233_out);

   SharedReg234_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_1_impl_out,
                 Y => SharedReg234_out);

   SharedReg235_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg234_out,
                 Y => SharedReg235_out);

   SharedReg236_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg235_out,
                 Y => SharedReg236_out);

   SharedReg237_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg236_out,
                 Y => SharedReg237_out);

   SharedReg238_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg237_out,
                 Y => SharedReg238_out);

   SharedReg239_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg238_out,
                 Y => SharedReg239_out);

   SharedReg240_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg239_out,
                 Y => SharedReg240_out);

   SharedReg241_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg240_out,
                 Y => SharedReg241_out);

   SharedReg242_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg241_out,
                 Y => SharedReg242_out);

   SharedReg243_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg242_out,
                 Y => SharedReg243_out);

   SharedReg244_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg243_out,
                 Y => SharedReg244_out);

   SharedReg245_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg244_out,
                 Y => SharedReg245_out);

   SharedReg246_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg245_out,
                 Y => SharedReg246_out);

   SharedReg247_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg246_out,
                 Y => SharedReg247_out);

   SharedReg248_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg247_out,
                 Y => SharedReg248_out);

   SharedReg249_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg248_out,
                 Y => SharedReg249_out);

   SharedReg250_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg249_out,
                 Y => SharedReg250_out);

   SharedReg251_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg250_out,
                 Y => SharedReg251_out);

   SharedReg252_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg251_out,
                 Y => SharedReg252_out);

   SharedReg253_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg252_out,
                 Y => SharedReg253_out);

   SharedReg254_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg253_out,
                 Y => SharedReg254_out);

   SharedReg255_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg254_out,
                 Y => SharedReg255_out);

   SharedReg256_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg255_out,
                 Y => SharedReg256_out);

   SharedReg257_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg256_out,
                 Y => SharedReg257_out);

   SharedReg258_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg257_out,
                 Y => SharedReg258_out);

   SharedReg259_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg258_out,
                 Y => SharedReg259_out);

   SharedReg260_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_2_impl_out,
                 Y => SharedReg260_out);

   SharedReg261_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg260_out,
                 Y => SharedReg261_out);

   SharedReg262_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg261_out,
                 Y => SharedReg262_out);

   SharedReg263_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg262_out,
                 Y => SharedReg263_out);

   SharedReg264_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg263_out,
                 Y => SharedReg264_out);

   SharedReg265_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg264_out,
                 Y => SharedReg265_out);

   SharedReg266_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg265_out,
                 Y => SharedReg266_out);

   SharedReg267_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg266_out,
                 Y => SharedReg267_out);

   SharedReg268_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg267_out,
                 Y => SharedReg268_out);

   SharedReg269_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg268_out,
                 Y => SharedReg269_out);

   SharedReg270_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg269_out,
                 Y => SharedReg270_out);

   SharedReg271_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg270_out,
                 Y => SharedReg271_out);

   SharedReg272_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg271_out,
                 Y => SharedReg272_out);

   SharedReg273_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg272_out,
                 Y => SharedReg273_out);

   SharedReg274_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg273_out,
                 Y => SharedReg274_out);

   SharedReg275_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg274_out,
                 Y => SharedReg275_out);

   SharedReg276_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg275_out,
                 Y => SharedReg276_out);

   SharedReg277_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg276_out,
                 Y => SharedReg277_out);

   SharedReg278_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg277_out,
                 Y => SharedReg278_out);

   SharedReg279_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg278_out,
                 Y => SharedReg279_out);

   SharedReg280_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg279_out,
                 Y => SharedReg280_out);

   SharedReg281_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg280_out,
                 Y => SharedReg281_out);

   SharedReg282_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg281_out,
                 Y => SharedReg282_out);

   SharedReg283_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg282_out,
                 Y => SharedReg283_out);

   SharedReg284_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg283_out,
                 Y => SharedReg284_out);

   SharedReg285_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_3_impl_out,
                 Y => SharedReg285_out);

   SharedReg286_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg285_out,
                 Y => SharedReg286_out);

   SharedReg287_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg286_out,
                 Y => SharedReg287_out);

   SharedReg288_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg287_out,
                 Y => SharedReg288_out);

   SharedReg289_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg288_out,
                 Y => SharedReg289_out);

   SharedReg290_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg289_out,
                 Y => SharedReg290_out);

   SharedReg291_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg290_out,
                 Y => SharedReg291_out);

   SharedReg292_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg291_out,
                 Y => SharedReg292_out);

   SharedReg293_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg292_out,
                 Y => SharedReg293_out);

   SharedReg294_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg293_out,
                 Y => SharedReg294_out);

   SharedReg295_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg294_out,
                 Y => SharedReg295_out);

   SharedReg296_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg295_out,
                 Y => SharedReg296_out);

   SharedReg297_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg296_out,
                 Y => SharedReg297_out);

   SharedReg298_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg297_out,
                 Y => SharedReg298_out);

   SharedReg299_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg298_out,
                 Y => SharedReg299_out);

   SharedReg300_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg299_out,
                 Y => SharedReg300_out);

   SharedReg301_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg300_out,
                 Y => SharedReg301_out);

   SharedReg302_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg301_out,
                 Y => SharedReg302_out);

   SharedReg303_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg302_out,
                 Y => SharedReg303_out);

   SharedReg304_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg303_out,
                 Y => SharedReg304_out);

   SharedReg305_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg304_out,
                 Y => SharedReg305_out);

   SharedReg306_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg305_out,
                 Y => SharedReg306_out);

   SharedReg307_instance: Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=30 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg306_out,
                 Y => SharedReg307_out);

   SharedReg308_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg307_out,
                 Y => SharedReg308_out);

   SharedReg309_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg308_out,
                 Y => SharedReg309_out);

   SharedReg310_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_4_impl_out,
                 Y => SharedReg310_out);

   SharedReg311_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg310_out,
                 Y => SharedReg311_out);

   SharedReg312_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg311_out,
                 Y => SharedReg312_out);

   SharedReg313_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg312_out,
                 Y => SharedReg313_out);

   SharedReg314_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg313_out,
                 Y => SharedReg314_out);

   SharedReg315_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg314_out,
                 Y => SharedReg315_out);

   SharedReg316_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg315_out,
                 Y => SharedReg316_out);

   SharedReg317_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg316_out,
                 Y => SharedReg317_out);

   SharedReg318_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg317_out,
                 Y => SharedReg318_out);

   SharedReg319_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg318_out,
                 Y => SharedReg319_out);

   SharedReg320_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg319_out,
                 Y => SharedReg320_out);

   SharedReg321_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg320_out,
                 Y => SharedReg321_out);

   SharedReg322_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg321_out,
                 Y => SharedReg322_out);

   SharedReg323_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg322_out,
                 Y => SharedReg323_out);

   SharedReg324_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg323_out,
                 Y => SharedReg324_out);

   SharedReg325_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg324_out,
                 Y => SharedReg325_out);

   SharedReg326_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg325_out,
                 Y => SharedReg326_out);

   SharedReg327_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg326_out,
                 Y => SharedReg327_out);

   SharedReg328_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg327_out,
                 Y => SharedReg328_out);

   SharedReg329_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg328_out,
                 Y => SharedReg329_out);

   SharedReg330_instance: Delay_34_DelayLength_38_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=38 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg329_out,
                 Y => SharedReg330_out);

   SharedReg331_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg330_out,
                 Y => SharedReg331_out);

   SharedReg332_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_6_impl_out,
                 Y => SharedReg332_out);

   SharedReg333_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg332_out,
                 Y => SharedReg333_out);

   SharedReg334_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg333_out,
                 Y => SharedReg334_out);

   SharedReg335_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg334_out,
                 Y => SharedReg335_out);

   SharedReg336_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg335_out,
                 Y => SharedReg336_out);

   SharedReg337_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg336_out,
                 Y => SharedReg337_out);

   SharedReg338_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg337_out,
                 Y => SharedReg338_out);

   SharedReg339_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg338_out,
                 Y => SharedReg339_out);

   SharedReg340_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg339_out,
                 Y => SharedReg340_out);

   SharedReg341_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg340_out,
                 Y => SharedReg341_out);

   SharedReg342_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg341_out,
                 Y => SharedReg342_out);

   SharedReg343_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg342_out,
                 Y => SharedReg343_out);

   SharedReg344_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg343_out,
                 Y => SharedReg344_out);

   SharedReg345_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg344_out,
                 Y => SharedReg345_out);

   SharedReg346_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg345_out,
                 Y => SharedReg346_out);

   SharedReg347_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg346_out,
                 Y => SharedReg347_out);

   SharedReg348_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg347_out,
                 Y => SharedReg348_out);

   SharedReg349_instance: Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=31 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg348_out,
                 Y => SharedReg349_out);

   SharedReg350_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_0_impl_out,
                 Y => SharedReg350_out);

   SharedReg351_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg350_out,
                 Y => SharedReg351_out);

   SharedReg352_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg351_out,
                 Y => SharedReg352_out);

   SharedReg353_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg352_out,
                 Y => SharedReg353_out);

   SharedReg354_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg353_out,
                 Y => SharedReg354_out);

   SharedReg355_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg354_out,
                 Y => SharedReg355_out);

   SharedReg356_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg355_out,
                 Y => SharedReg356_out);

   SharedReg357_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg356_out,
                 Y => SharedReg357_out);

   SharedReg358_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg357_out,
                 Y => SharedReg358_out);

   SharedReg359_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg358_out,
                 Y => SharedReg359_out);

   SharedReg360_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg359_out,
                 Y => SharedReg360_out);

   SharedReg361_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg360_out,
                 Y => SharedReg361_out);

   SharedReg362_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg361_out,
                 Y => SharedReg362_out);

   SharedReg363_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg362_out,
                 Y => SharedReg363_out);

   SharedReg364_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg363_out,
                 Y => SharedReg364_out);

   SharedReg365_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_1_impl_out,
                 Y => SharedReg365_out);

   SharedReg366_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg365_out,
                 Y => SharedReg366_out);

   SharedReg367_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg366_out,
                 Y => SharedReg367_out);

   SharedReg368_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg367_out,
                 Y => SharedReg368_out);

   SharedReg369_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg368_out,
                 Y => SharedReg369_out);

   SharedReg370_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg369_out,
                 Y => SharedReg370_out);

   SharedReg371_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg370_out,
                 Y => SharedReg371_out);

   SharedReg372_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg371_out,
                 Y => SharedReg372_out);

   SharedReg373_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg372_out,
                 Y => SharedReg373_out);

   SharedReg374_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg373_out,
                 Y => SharedReg374_out);

   SharedReg375_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg374_out,
                 Y => SharedReg375_out);

   SharedReg376_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg375_out,
                 Y => SharedReg376_out);

   SharedReg377_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg376_out,
                 Y => SharedReg377_out);

   SharedReg378_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg377_out,
                 Y => SharedReg378_out);

   SharedReg379_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg378_out,
                 Y => SharedReg379_out);

   SharedReg380_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_2_impl_out,
                 Y => SharedReg380_out);

   SharedReg381_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg380_out,
                 Y => SharedReg381_out);

   SharedReg382_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg381_out,
                 Y => SharedReg382_out);

   SharedReg383_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg382_out,
                 Y => SharedReg383_out);

   SharedReg384_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg383_out,
                 Y => SharedReg384_out);

   SharedReg385_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg384_out,
                 Y => SharedReg385_out);

   SharedReg386_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg385_out,
                 Y => SharedReg386_out);

   SharedReg387_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg386_out,
                 Y => SharedReg387_out);

   SharedReg388_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg387_out,
                 Y => SharedReg388_out);

   SharedReg389_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg388_out,
                 Y => SharedReg389_out);

   SharedReg390_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg389_out,
                 Y => SharedReg390_out);

   SharedReg391_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg390_out,
                 Y => SharedReg391_out);

   SharedReg392_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg391_out,
                 Y => SharedReg392_out);

   SharedReg393_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg392_out,
                 Y => SharedReg393_out);

   SharedReg394_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg393_out,
                 Y => SharedReg394_out);

   SharedReg395_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_3_impl_out,
                 Y => SharedReg395_out);

   SharedReg396_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg395_out,
                 Y => SharedReg396_out);

   SharedReg397_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg396_out,
                 Y => SharedReg397_out);

   SharedReg398_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg397_out,
                 Y => SharedReg398_out);

   SharedReg399_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg398_out,
                 Y => SharedReg399_out);

   SharedReg400_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg399_out,
                 Y => SharedReg400_out);

   SharedReg401_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg400_out,
                 Y => SharedReg401_out);

   SharedReg402_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg401_out,
                 Y => SharedReg402_out);

   SharedReg403_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg402_out,
                 Y => SharedReg403_out);

   SharedReg404_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg403_out,
                 Y => SharedReg404_out);

   SharedReg405_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg404_out,
                 Y => SharedReg405_out);

   SharedReg406_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg405_out,
                 Y => SharedReg406_out);

   SharedReg407_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg406_out,
                 Y => SharedReg407_out);

   SharedReg408_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg407_out,
                 Y => SharedReg408_out);

   SharedReg409_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg408_out,
                 Y => SharedReg409_out);

   SharedReg410_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_4_impl_out,
                 Y => SharedReg410_out);

   SharedReg411_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg410_out,
                 Y => SharedReg411_out);

   SharedReg412_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg411_out,
                 Y => SharedReg412_out);

   SharedReg413_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg412_out,
                 Y => SharedReg413_out);

   SharedReg414_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg413_out,
                 Y => SharedReg414_out);

   SharedReg415_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg414_out,
                 Y => SharedReg415_out);

   SharedReg416_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg415_out,
                 Y => SharedReg416_out);

   SharedReg417_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg416_out,
                 Y => SharedReg417_out);

   SharedReg418_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg417_out,
                 Y => SharedReg418_out);

   SharedReg419_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg418_out,
                 Y => SharedReg419_out);

   SharedReg420_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg419_out,
                 Y => SharedReg420_out);

   SharedReg421_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg420_out,
                 Y => SharedReg421_out);

   SharedReg422_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg421_out,
                 Y => SharedReg422_out);

   SharedReg423_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg422_out,
                 Y => SharedReg423_out);

   SharedReg424_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg423_out,
                 Y => SharedReg424_out);

   SharedReg425_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_5_impl_out,
                 Y => SharedReg425_out);

   SharedReg426_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg425_out,
                 Y => SharedReg426_out);

   SharedReg427_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg426_out,
                 Y => SharedReg427_out);

   SharedReg428_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg427_out,
                 Y => SharedReg428_out);

   SharedReg429_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg428_out,
                 Y => SharedReg429_out);

   SharedReg430_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg429_out,
                 Y => SharedReg430_out);

   SharedReg431_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg430_out,
                 Y => SharedReg431_out);

   SharedReg432_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg431_out,
                 Y => SharedReg432_out);

   SharedReg433_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg432_out,
                 Y => SharedReg433_out);

   SharedReg434_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg433_out,
                 Y => SharedReg434_out);

   SharedReg435_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg434_out,
                 Y => SharedReg435_out);

   SharedReg436_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg435_out,
                 Y => SharedReg436_out);

   SharedReg437_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg436_out,
                 Y => SharedReg437_out);

   SharedReg438_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg437_out,
                 Y => SharedReg438_out);

   SharedReg439_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg438_out,
                 Y => SharedReg439_out);

   SharedReg440_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_6_impl_out,
                 Y => SharedReg440_out);

   SharedReg441_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg440_out,
                 Y => SharedReg441_out);

   SharedReg442_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg441_out,
                 Y => SharedReg442_out);

   SharedReg443_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg442_out,
                 Y => SharedReg443_out);

   SharedReg444_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg443_out,
                 Y => SharedReg444_out);

   SharedReg445_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg444_out,
                 Y => SharedReg445_out);

   SharedReg446_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg445_out,
                 Y => SharedReg446_out);

   SharedReg447_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg446_out,
                 Y => SharedReg447_out);

   SharedReg448_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg447_out,
                 Y => SharedReg448_out);

   SharedReg449_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg448_out,
                 Y => SharedReg449_out);

   SharedReg450_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg449_out,
                 Y => SharedReg450_out);

   SharedReg451_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg450_out,
                 Y => SharedReg451_out);

   SharedReg452_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg451_out,
                 Y => SharedReg452_out);

   SharedReg453_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg452_out,
                 Y => SharedReg453_out);

   SharedReg454_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg453_out,
                 Y => SharedReg454_out);

   SharedReg455_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product31_0_impl_out,
                 Y => SharedReg455_out);

   SharedReg456_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg455_out,
                 Y => SharedReg456_out);

   SharedReg457_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg456_out,
                 Y => SharedReg457_out);

   SharedReg458_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg457_out,
                 Y => SharedReg458_out);

   SharedReg459_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg458_out,
                 Y => SharedReg459_out);

   SharedReg460_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg459_out,
                 Y => SharedReg460_out);

   SharedReg461_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg460_out,
                 Y => SharedReg461_out);

   SharedReg462_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg461_out,
                 Y => SharedReg462_out);

   SharedReg463_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg462_out,
                 Y => SharedReg463_out);

   SharedReg464_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg463_out,
                 Y => SharedReg464_out);

   SharedReg465_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg464_out,
                 Y => SharedReg465_out);

   SharedReg466_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg465_out,
                 Y => SharedReg466_out);

   SharedReg467_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg466_out,
                 Y => SharedReg467_out);

   SharedReg468_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg467_out,
                 Y => SharedReg468_out);

   SharedReg469_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg468_out,
                 Y => SharedReg469_out);

   SharedReg470_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg469_out,
                 Y => SharedReg470_out);

   SharedReg471_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product31_1_impl_out,
                 Y => SharedReg471_out);

   SharedReg472_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg471_out,
                 Y => SharedReg472_out);

   SharedReg473_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg472_out,
                 Y => SharedReg473_out);

   SharedReg474_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg473_out,
                 Y => SharedReg474_out);

   SharedReg475_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg474_out,
                 Y => SharedReg475_out);

   SharedReg476_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg475_out,
                 Y => SharedReg476_out);

   SharedReg477_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg476_out,
                 Y => SharedReg477_out);

   SharedReg478_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg477_out,
                 Y => SharedReg478_out);

   SharedReg479_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg478_out,
                 Y => SharedReg479_out);

   SharedReg480_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg479_out,
                 Y => SharedReg480_out);

   SharedReg481_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg480_out,
                 Y => SharedReg481_out);

   SharedReg482_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg481_out,
                 Y => SharedReg482_out);

   SharedReg483_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg482_out,
                 Y => SharedReg483_out);

   SharedReg484_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg483_out,
                 Y => SharedReg484_out);

   SharedReg485_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg484_out,
                 Y => SharedReg485_out);

   SharedReg486_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg485_out,
                 Y => SharedReg486_out);

   SharedReg487_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product31_2_impl_out,
                 Y => SharedReg487_out);

   SharedReg488_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg487_out,
                 Y => SharedReg488_out);

   SharedReg489_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg488_out,
                 Y => SharedReg489_out);

   SharedReg490_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg489_out,
                 Y => SharedReg490_out);

   SharedReg491_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg490_out,
                 Y => SharedReg491_out);

   SharedReg492_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg491_out,
                 Y => SharedReg492_out);

   SharedReg493_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg492_out,
                 Y => SharedReg493_out);

   SharedReg494_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg493_out,
                 Y => SharedReg494_out);

   SharedReg495_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg494_out,
                 Y => SharedReg495_out);

   SharedReg496_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg495_out,
                 Y => SharedReg496_out);

   SharedReg497_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg496_out,
                 Y => SharedReg497_out);

   SharedReg498_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg497_out,
                 Y => SharedReg498_out);

   SharedReg499_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg498_out,
                 Y => SharedReg499_out);

   SharedReg500_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg499_out,
                 Y => SharedReg500_out);

   SharedReg501_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg500_out,
                 Y => SharedReg501_out);

   SharedReg502_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg501_out,
                 Y => SharedReg502_out);

   SharedReg503_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product31_3_impl_out,
                 Y => SharedReg503_out);

   SharedReg504_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg503_out,
                 Y => SharedReg504_out);

   SharedReg505_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg504_out,
                 Y => SharedReg505_out);

   SharedReg506_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg505_out,
                 Y => SharedReg506_out);

   SharedReg507_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg506_out,
                 Y => SharedReg507_out);

   SharedReg508_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg507_out,
                 Y => SharedReg508_out);

   SharedReg509_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg508_out,
                 Y => SharedReg509_out);

   SharedReg510_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg509_out,
                 Y => SharedReg510_out);

   SharedReg511_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg510_out,
                 Y => SharedReg511_out);

   SharedReg512_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg511_out,
                 Y => SharedReg512_out);

   SharedReg513_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg512_out,
                 Y => SharedReg513_out);

   SharedReg514_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg513_out,
                 Y => SharedReg514_out);

   SharedReg515_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg514_out,
                 Y => SharedReg515_out);

   SharedReg516_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg515_out,
                 Y => SharedReg516_out);

   SharedReg517_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg516_out,
                 Y => SharedReg517_out);

   SharedReg518_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg517_out,
                 Y => SharedReg518_out);

   SharedReg519_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product31_4_impl_out,
                 Y => SharedReg519_out);

   SharedReg520_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg519_out,
                 Y => SharedReg520_out);

   SharedReg521_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg520_out,
                 Y => SharedReg521_out);

   SharedReg522_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg521_out,
                 Y => SharedReg522_out);

   SharedReg523_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg522_out,
                 Y => SharedReg523_out);

   SharedReg524_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg523_out,
                 Y => SharedReg524_out);

   SharedReg525_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg524_out,
                 Y => SharedReg525_out);

   SharedReg526_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg525_out,
                 Y => SharedReg526_out);

   SharedReg527_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg526_out,
                 Y => SharedReg527_out);

   SharedReg528_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg527_out,
                 Y => SharedReg528_out);

   SharedReg529_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg528_out,
                 Y => SharedReg529_out);

   SharedReg530_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg529_out,
                 Y => SharedReg530_out);

   SharedReg531_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg530_out,
                 Y => SharedReg531_out);

   SharedReg532_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg531_out,
                 Y => SharedReg532_out);

   SharedReg533_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg532_out,
                 Y => SharedReg533_out);

   SharedReg534_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg533_out,
                 Y => SharedReg534_out);

   SharedReg535_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product31_5_impl_out,
                 Y => SharedReg535_out);

   SharedReg536_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg535_out,
                 Y => SharedReg536_out);

   SharedReg537_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg536_out,
                 Y => SharedReg537_out);

   SharedReg538_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg537_out,
                 Y => SharedReg538_out);

   SharedReg539_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg538_out,
                 Y => SharedReg539_out);

   SharedReg540_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg539_out,
                 Y => SharedReg540_out);

   SharedReg541_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg540_out,
                 Y => SharedReg541_out);

   SharedReg542_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg541_out,
                 Y => SharedReg542_out);

   SharedReg543_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg542_out,
                 Y => SharedReg543_out);

   SharedReg544_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg543_out,
                 Y => SharedReg544_out);

   SharedReg545_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg544_out,
                 Y => SharedReg545_out);

   SharedReg546_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg545_out,
                 Y => SharedReg546_out);

   SharedReg547_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg546_out,
                 Y => SharedReg547_out);

   SharedReg548_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg547_out,
                 Y => SharedReg548_out);

   SharedReg549_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg548_out,
                 Y => SharedReg549_out);

   SharedReg550_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg549_out,
                 Y => SharedReg550_out);

   SharedReg551_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product31_6_impl_out,
                 Y => SharedReg551_out);

   SharedReg552_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg551_out,
                 Y => SharedReg552_out);

   SharedReg553_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg552_out,
                 Y => SharedReg553_out);

   SharedReg554_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg553_out,
                 Y => SharedReg554_out);

   SharedReg555_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg554_out,
                 Y => SharedReg555_out);

   SharedReg556_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg555_out,
                 Y => SharedReg556_out);

   SharedReg557_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg556_out,
                 Y => SharedReg557_out);

   SharedReg558_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg557_out,
                 Y => SharedReg558_out);

   SharedReg559_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg558_out,
                 Y => SharedReg559_out);

   SharedReg560_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg559_out,
                 Y => SharedReg560_out);

   SharedReg561_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg560_out,
                 Y => SharedReg561_out);

   SharedReg562_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg561_out,
                 Y => SharedReg562_out);

   SharedReg563_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg562_out,
                 Y => SharedReg563_out);

   SharedReg564_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg563_out,
                 Y => SharedReg564_out);

   SharedReg565_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg564_out,
                 Y => SharedReg565_out);

   SharedReg566_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg565_out,
                 Y => SharedReg566_out);

   SharedReg567_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_0_impl_out,
                 Y => SharedReg567_out);

   SharedReg568_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg567_out,
                 Y => SharedReg568_out);

   SharedReg569_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg568_out,
                 Y => SharedReg569_out);

   SharedReg570_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg569_out,
                 Y => SharedReg570_out);

   SharedReg571_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg570_out,
                 Y => SharedReg571_out);

   SharedReg572_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg571_out,
                 Y => SharedReg572_out);

   SharedReg573_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg572_out,
                 Y => SharedReg573_out);

   SharedReg574_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg573_out,
                 Y => SharedReg574_out);

   SharedReg575_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg574_out,
                 Y => SharedReg575_out);

   SharedReg576_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg575_out,
                 Y => SharedReg576_out);

   SharedReg577_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg576_out,
                 Y => SharedReg577_out);

   SharedReg578_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg577_out,
                 Y => SharedReg578_out);

   SharedReg579_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg578_out,
                 Y => SharedReg579_out);

   SharedReg580_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg579_out,
                 Y => SharedReg580_out);

   SharedReg581_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg580_out,
                 Y => SharedReg581_out);

   SharedReg582_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg581_out,
                 Y => SharedReg582_out);

   SharedReg583_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg582_out,
                 Y => SharedReg583_out);

   SharedReg584_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg583_out,
                 Y => SharedReg584_out);

   SharedReg585_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg584_out,
                 Y => SharedReg585_out);

   SharedReg586_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg585_out,
                 Y => SharedReg586_out);

   SharedReg587_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg586_out,
                 Y => SharedReg587_out);

   SharedReg588_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg587_out,
                 Y => SharedReg588_out);

   SharedReg589_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg588_out,
                 Y => SharedReg589_out);

   SharedReg590_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg589_out,
                 Y => SharedReg590_out);

   SharedReg591_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg590_out,
                 Y => SharedReg591_out);

   SharedReg592_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg591_out,
                 Y => SharedReg592_out);

   SharedReg593_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_1_impl_out,
                 Y => SharedReg593_out);

   SharedReg594_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg593_out,
                 Y => SharedReg594_out);

   SharedReg595_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg594_out,
                 Y => SharedReg595_out);

   SharedReg596_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg595_out,
                 Y => SharedReg596_out);

   SharedReg597_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg596_out,
                 Y => SharedReg597_out);

   SharedReg598_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg597_out,
                 Y => SharedReg598_out);

   SharedReg599_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg598_out,
                 Y => SharedReg599_out);

   SharedReg600_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg599_out,
                 Y => SharedReg600_out);

   SharedReg601_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg600_out,
                 Y => SharedReg601_out);

   SharedReg602_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg601_out,
                 Y => SharedReg602_out);

   SharedReg603_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg602_out,
                 Y => SharedReg603_out);

   SharedReg604_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg603_out,
                 Y => SharedReg604_out);

   SharedReg605_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg604_out,
                 Y => SharedReg605_out);

   SharedReg606_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg605_out,
                 Y => SharedReg606_out);

   SharedReg607_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg606_out,
                 Y => SharedReg607_out);

   SharedReg608_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg607_out,
                 Y => SharedReg608_out);

   SharedReg609_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg608_out,
                 Y => SharedReg609_out);

   SharedReg610_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg609_out,
                 Y => SharedReg610_out);

   SharedReg611_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg610_out,
                 Y => SharedReg611_out);

   SharedReg612_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg611_out,
                 Y => SharedReg612_out);

   SharedReg613_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg612_out,
                 Y => SharedReg613_out);

   SharedReg614_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg613_out,
                 Y => SharedReg614_out);

   SharedReg615_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg614_out,
                 Y => SharedReg615_out);

   SharedReg616_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg615_out,
                 Y => SharedReg616_out);

   SharedReg617_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_2_impl_out,
                 Y => SharedReg617_out);

   SharedReg618_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg617_out,
                 Y => SharedReg618_out);

   SharedReg619_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg618_out,
                 Y => SharedReg619_out);

   SharedReg620_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg619_out,
                 Y => SharedReg620_out);

   SharedReg621_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg620_out,
                 Y => SharedReg621_out);

   SharedReg622_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg621_out,
                 Y => SharedReg622_out);

   SharedReg623_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg622_out,
                 Y => SharedReg623_out);

   SharedReg624_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg623_out,
                 Y => SharedReg624_out);

   SharedReg625_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg624_out,
                 Y => SharedReg625_out);

   SharedReg626_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg625_out,
                 Y => SharedReg626_out);

   SharedReg627_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg626_out,
                 Y => SharedReg627_out);

   SharedReg628_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg627_out,
                 Y => SharedReg628_out);

   SharedReg629_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg628_out,
                 Y => SharedReg629_out);

   SharedReg630_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg629_out,
                 Y => SharedReg630_out);

   SharedReg631_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg630_out,
                 Y => SharedReg631_out);

   SharedReg632_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg631_out,
                 Y => SharedReg632_out);

   SharedReg633_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg632_out,
                 Y => SharedReg633_out);

   SharedReg634_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg633_out,
                 Y => SharedReg634_out);

   SharedReg635_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg634_out,
                 Y => SharedReg635_out);

   SharedReg636_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg635_out,
                 Y => SharedReg636_out);

   SharedReg637_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg636_out,
                 Y => SharedReg637_out);

   SharedReg638_instance: Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=30 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg637_out,
                 Y => SharedReg638_out);

   SharedReg639_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg638_out,
                 Y => SharedReg639_out);

   SharedReg640_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_3_impl_out,
                 Y => SharedReg640_out);

   SharedReg641_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg640_out,
                 Y => SharedReg641_out);

   SharedReg642_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg641_out,
                 Y => SharedReg642_out);

   SharedReg643_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg642_out,
                 Y => SharedReg643_out);

   SharedReg644_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg643_out,
                 Y => SharedReg644_out);

   SharedReg645_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg644_out,
                 Y => SharedReg645_out);

   SharedReg646_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg645_out,
                 Y => SharedReg646_out);

   SharedReg647_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg646_out,
                 Y => SharedReg647_out);

   SharedReg648_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg647_out,
                 Y => SharedReg648_out);

   SharedReg649_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg648_out,
                 Y => SharedReg649_out);

   SharedReg650_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg649_out,
                 Y => SharedReg650_out);

   SharedReg651_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg650_out,
                 Y => SharedReg651_out);

   SharedReg652_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg651_out,
                 Y => SharedReg652_out);

   SharedReg653_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg652_out,
                 Y => SharedReg653_out);

   SharedReg654_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg653_out,
                 Y => SharedReg654_out);

   SharedReg655_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg654_out,
                 Y => SharedReg655_out);

   SharedReg656_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg655_out,
                 Y => SharedReg656_out);

   SharedReg657_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg656_out,
                 Y => SharedReg657_out);

   SharedReg658_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg657_out,
                 Y => SharedReg658_out);

   SharedReg659_instance: Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=30 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg658_out,
                 Y => SharedReg659_out);

   SharedReg660_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg659_out,
                 Y => SharedReg660_out);

   SharedReg661_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_4_impl_out,
                 Y => SharedReg661_out);

   SharedReg662_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg661_out,
                 Y => SharedReg662_out);

   SharedReg663_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg662_out,
                 Y => SharedReg663_out);

   SharedReg664_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg663_out,
                 Y => SharedReg664_out);

   SharedReg665_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg664_out,
                 Y => SharedReg665_out);

   SharedReg666_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg665_out,
                 Y => SharedReg666_out);

   SharedReg667_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg666_out,
                 Y => SharedReg667_out);

   SharedReg668_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg667_out,
                 Y => SharedReg668_out);

   SharedReg669_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg668_out,
                 Y => SharedReg669_out);

   SharedReg670_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg669_out,
                 Y => SharedReg670_out);

   SharedReg671_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg670_out,
                 Y => SharedReg671_out);

   SharedReg672_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg671_out,
                 Y => SharedReg672_out);

   SharedReg673_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg672_out,
                 Y => SharedReg673_out);

   SharedReg674_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg673_out,
                 Y => SharedReg674_out);

   SharedReg675_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg674_out,
                 Y => SharedReg675_out);

   SharedReg676_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg675_out,
                 Y => SharedReg676_out);

   SharedReg677_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg676_out,
                 Y => SharedReg677_out);

   SharedReg678_instance: Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=22 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg677_out,
                 Y => SharedReg678_out);

   SharedReg679_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg678_out,
                 Y => SharedReg679_out);

   SharedReg680_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg679_out,
                 Y => SharedReg680_out);

   SharedReg681_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg680_out,
                 Y => SharedReg681_out);

   SharedReg682_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg681_out,
                 Y => SharedReg682_out);

   SharedReg683_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg682_out,
                 Y => SharedReg683_out);

   SharedReg684_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg683_out,
                 Y => SharedReg684_out);

   SharedReg685_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_5_impl_out,
                 Y => SharedReg685_out);

   SharedReg686_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg685_out,
                 Y => SharedReg686_out);

   SharedReg687_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg686_out,
                 Y => SharedReg687_out);

   SharedReg688_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg687_out,
                 Y => SharedReg688_out);

   SharedReg689_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg688_out,
                 Y => SharedReg689_out);

   SharedReg690_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg689_out,
                 Y => SharedReg690_out);

   SharedReg691_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg690_out,
                 Y => SharedReg691_out);

   SharedReg692_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg691_out,
                 Y => SharedReg692_out);

   SharedReg693_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg692_out,
                 Y => SharedReg693_out);

   SharedReg694_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg693_out,
                 Y => SharedReg694_out);

   SharedReg695_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg694_out,
                 Y => SharedReg695_out);

   SharedReg696_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg695_out,
                 Y => SharedReg696_out);

   SharedReg697_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg696_out,
                 Y => SharedReg697_out);

   SharedReg698_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg697_out,
                 Y => SharedReg698_out);

   SharedReg699_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg698_out,
                 Y => SharedReg699_out);

   SharedReg700_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg699_out,
                 Y => SharedReg700_out);

   SharedReg701_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg700_out,
                 Y => SharedReg701_out);

   SharedReg702_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg701_out,
                 Y => SharedReg702_out);

   SharedReg703_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg702_out,
                 Y => SharedReg703_out);

   SharedReg704_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg703_out,
                 Y => SharedReg704_out);

   SharedReg705_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg704_out,
                 Y => SharedReg705_out);

   SharedReg706_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg705_out,
                 Y => SharedReg706_out);

   SharedReg707_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_6_impl_out,
                 Y => SharedReg707_out);

   SharedReg708_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg707_out,
                 Y => SharedReg708_out);

   SharedReg709_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg708_out,
                 Y => SharedReg709_out);

   SharedReg710_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg709_out,
                 Y => SharedReg710_out);

   SharedReg711_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg710_out,
                 Y => SharedReg711_out);

   SharedReg712_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg711_out,
                 Y => SharedReg712_out);

   SharedReg713_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg712_out,
                 Y => SharedReg713_out);

   SharedReg714_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg713_out,
                 Y => SharedReg714_out);

   SharedReg715_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg714_out,
                 Y => SharedReg715_out);

   SharedReg716_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg715_out,
                 Y => SharedReg716_out);

   SharedReg717_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg716_out,
                 Y => SharedReg717_out);

   SharedReg718_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg717_out,
                 Y => SharedReg718_out);

   SharedReg719_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg718_out,
                 Y => SharedReg719_out);

   SharedReg720_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg719_out,
                 Y => SharedReg720_out);

   SharedReg721_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg720_out,
                 Y => SharedReg721_out);

   SharedReg722_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg721_out,
                 Y => SharedReg722_out);

   SharedReg723_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg722_out,
                 Y => SharedReg723_out);

   SharedReg724_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg723_out,
                 Y => SharedReg724_out);

   SharedReg725_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg724_out,
                 Y => SharedReg725_out);

   SharedReg726_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg725_out,
                 Y => SharedReg726_out);

   SharedReg727_instance: Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=28 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg726_out,
                 Y => SharedReg727_out);

   SharedReg728_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg727_out,
                 Y => SharedReg728_out);

   SharedReg729_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_0_impl_out,
                 Y => SharedReg729_out);

   SharedReg730_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg729_out,
                 Y => SharedReg730_out);

   SharedReg731_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg730_out,
                 Y => SharedReg731_out);

   SharedReg732_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg731_out,
                 Y => SharedReg732_out);

   SharedReg733_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg732_out,
                 Y => SharedReg733_out);

   SharedReg734_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg733_out,
                 Y => SharedReg734_out);

   SharedReg735_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg734_out,
                 Y => SharedReg735_out);

   SharedReg736_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg735_out,
                 Y => SharedReg736_out);

   SharedReg737_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg736_out,
                 Y => SharedReg737_out);

   SharedReg738_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg737_out,
                 Y => SharedReg738_out);

   SharedReg739_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg738_out,
                 Y => SharedReg739_out);

   SharedReg740_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg739_out,
                 Y => SharedReg740_out);

   SharedReg741_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg740_out,
                 Y => SharedReg741_out);

   SharedReg742_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg741_out,
                 Y => SharedReg742_out);

   SharedReg743_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg742_out,
                 Y => SharedReg743_out);

   SharedReg744_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg743_out,
                 Y => SharedReg744_out);

   SharedReg745_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg744_out,
                 Y => SharedReg745_out);

   SharedReg746_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg745_out,
                 Y => SharedReg746_out);

   SharedReg747_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_1_impl_out,
                 Y => SharedReg747_out);

   SharedReg748_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg747_out,
                 Y => SharedReg748_out);

   SharedReg749_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg748_out,
                 Y => SharedReg749_out);

   SharedReg750_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg749_out,
                 Y => SharedReg750_out);

   SharedReg751_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg750_out,
                 Y => SharedReg751_out);

   SharedReg752_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg751_out,
                 Y => SharedReg752_out);

   SharedReg753_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg752_out,
                 Y => SharedReg753_out);

   SharedReg754_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg753_out,
                 Y => SharedReg754_out);

   SharedReg755_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg754_out,
                 Y => SharedReg755_out);

   SharedReg756_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg755_out,
                 Y => SharedReg756_out);

   SharedReg757_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg756_out,
                 Y => SharedReg757_out);

   SharedReg758_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg757_out,
                 Y => SharedReg758_out);

   SharedReg759_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg758_out,
                 Y => SharedReg759_out);

   SharedReg760_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg759_out,
                 Y => SharedReg760_out);

   SharedReg761_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg760_out,
                 Y => SharedReg761_out);

   SharedReg762_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg761_out,
                 Y => SharedReg762_out);

   SharedReg763_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg762_out,
                 Y => SharedReg763_out);

   SharedReg764_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg763_out,
                 Y => SharedReg764_out);

   SharedReg765_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_2_impl_out,
                 Y => SharedReg765_out);

   SharedReg766_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg765_out,
                 Y => SharedReg766_out);

   SharedReg767_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg766_out,
                 Y => SharedReg767_out);

   SharedReg768_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg767_out,
                 Y => SharedReg768_out);

   SharedReg769_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg768_out,
                 Y => SharedReg769_out);

   SharedReg770_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg769_out,
                 Y => SharedReg770_out);

   SharedReg771_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg770_out,
                 Y => SharedReg771_out);

   SharedReg772_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg771_out,
                 Y => SharedReg772_out);

   SharedReg773_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg772_out,
                 Y => SharedReg773_out);

   SharedReg774_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg773_out,
                 Y => SharedReg774_out);

   SharedReg775_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg774_out,
                 Y => SharedReg775_out);

   SharedReg776_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg775_out,
                 Y => SharedReg776_out);

   SharedReg777_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg776_out,
                 Y => SharedReg777_out);

   SharedReg778_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg777_out,
                 Y => SharedReg778_out);

   SharedReg779_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg778_out,
                 Y => SharedReg779_out);

   SharedReg780_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg779_out,
                 Y => SharedReg780_out);

   SharedReg781_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg780_out,
                 Y => SharedReg781_out);

   SharedReg782_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg781_out,
                 Y => SharedReg782_out);

   SharedReg783_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_3_impl_out,
                 Y => SharedReg783_out);

   SharedReg784_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg783_out,
                 Y => SharedReg784_out);

   SharedReg785_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg784_out,
                 Y => SharedReg785_out);

   SharedReg786_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg785_out,
                 Y => SharedReg786_out);

   SharedReg787_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg786_out,
                 Y => SharedReg787_out);

   SharedReg788_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg787_out,
                 Y => SharedReg788_out);

   SharedReg789_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg788_out,
                 Y => SharedReg789_out);

   SharedReg790_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg789_out,
                 Y => SharedReg790_out);

   SharedReg791_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg790_out,
                 Y => SharedReg791_out);

   SharedReg792_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg791_out,
                 Y => SharedReg792_out);

   SharedReg793_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg792_out,
                 Y => SharedReg793_out);

   SharedReg794_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg793_out,
                 Y => SharedReg794_out);

   SharedReg795_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg794_out,
                 Y => SharedReg795_out);

   SharedReg796_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg795_out,
                 Y => SharedReg796_out);

   SharedReg797_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg796_out,
                 Y => SharedReg797_out);

   SharedReg798_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg797_out,
                 Y => SharedReg798_out);

   SharedReg799_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg798_out,
                 Y => SharedReg799_out);

   SharedReg800_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg799_out,
                 Y => SharedReg800_out);

   SharedReg801_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_4_impl_out,
                 Y => SharedReg801_out);

   SharedReg802_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg801_out,
                 Y => SharedReg802_out);

   SharedReg803_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg802_out,
                 Y => SharedReg803_out);

   SharedReg804_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg803_out,
                 Y => SharedReg804_out);

   SharedReg805_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg804_out,
                 Y => SharedReg805_out);

   SharedReg806_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg805_out,
                 Y => SharedReg806_out);

   SharedReg807_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg806_out,
                 Y => SharedReg807_out);

   SharedReg808_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg807_out,
                 Y => SharedReg808_out);

   SharedReg809_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg808_out,
                 Y => SharedReg809_out);

   SharedReg810_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg809_out,
                 Y => SharedReg810_out);

   SharedReg811_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg810_out,
                 Y => SharedReg811_out);

   SharedReg812_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg811_out,
                 Y => SharedReg812_out);

   SharedReg813_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg812_out,
                 Y => SharedReg813_out);

   SharedReg814_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg813_out,
                 Y => SharedReg814_out);

   SharedReg815_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg814_out,
                 Y => SharedReg815_out);

   SharedReg816_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg815_out,
                 Y => SharedReg816_out);

   SharedReg817_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg816_out,
                 Y => SharedReg817_out);

   SharedReg818_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg817_out,
                 Y => SharedReg818_out);

   SharedReg819_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_5_impl_out,
                 Y => SharedReg819_out);

   SharedReg820_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg819_out,
                 Y => SharedReg820_out);

   SharedReg821_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg820_out,
                 Y => SharedReg821_out);

   SharedReg822_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg821_out,
                 Y => SharedReg822_out);

   SharedReg823_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg822_out,
                 Y => SharedReg823_out);

   SharedReg824_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg823_out,
                 Y => SharedReg824_out);

   SharedReg825_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg824_out,
                 Y => SharedReg825_out);

   SharedReg826_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg825_out,
                 Y => SharedReg826_out);

   SharedReg827_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg826_out,
                 Y => SharedReg827_out);

   SharedReg828_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg827_out,
                 Y => SharedReg828_out);

   SharedReg829_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg828_out,
                 Y => SharedReg829_out);

   SharedReg830_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg829_out,
                 Y => SharedReg830_out);

   SharedReg831_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg830_out,
                 Y => SharedReg831_out);

   SharedReg832_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg831_out,
                 Y => SharedReg832_out);

   SharedReg833_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg832_out,
                 Y => SharedReg833_out);

   SharedReg834_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg833_out,
                 Y => SharedReg834_out);

   SharedReg835_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg834_out,
                 Y => SharedReg835_out);

   SharedReg836_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg835_out,
                 Y => SharedReg836_out);

   SharedReg837_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_6_impl_out,
                 Y => SharedReg837_out);

   SharedReg838_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg837_out,
                 Y => SharedReg838_out);

   SharedReg839_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg838_out,
                 Y => SharedReg839_out);

   SharedReg840_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg839_out,
                 Y => SharedReg840_out);

   SharedReg841_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg840_out,
                 Y => SharedReg841_out);

   SharedReg842_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg841_out,
                 Y => SharedReg842_out);

   SharedReg843_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg842_out,
                 Y => SharedReg843_out);

   SharedReg844_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg843_out,
                 Y => SharedReg844_out);

   SharedReg845_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg844_out,
                 Y => SharedReg845_out);

   SharedReg846_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg845_out,
                 Y => SharedReg846_out);

   SharedReg847_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg846_out,
                 Y => SharedReg847_out);

   SharedReg848_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg847_out,
                 Y => SharedReg848_out);

   SharedReg849_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg848_out,
                 Y => SharedReg849_out);

   SharedReg850_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg849_out,
                 Y => SharedReg850_out);

   SharedReg851_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg850_out,
                 Y => SharedReg851_out);

   SharedReg852_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg851_out,
                 Y => SharedReg852_out);

   SharedReg853_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg852_out,
                 Y => SharedReg853_out);

   SharedReg854_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg853_out,
                 Y => SharedReg854_out);

   SharedReg855_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract3_4_impl_out,
                 Y => SharedReg855_out);

   SharedReg856_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg855_out,
                 Y => SharedReg856_out);

   SharedReg857_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg856_out,
                 Y => SharedReg857_out);

   SharedReg858_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg857_out,
                 Y => SharedReg858_out);

   SharedReg859_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg858_out,
                 Y => SharedReg859_out);

   SharedReg860_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg859_out,
                 Y => SharedReg860_out);

   SharedReg861_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg860_out,
                 Y => SharedReg861_out);

   SharedReg862_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg861_out,
                 Y => SharedReg862_out);

   SharedReg863_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg862_out,
                 Y => SharedReg863_out);

   SharedReg864_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg863_out,
                 Y => SharedReg864_out);

   SharedReg865_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg864_out,
                 Y => SharedReg865_out);

   SharedReg866_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg865_out,
                 Y => SharedReg866_out);

   SharedReg867_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg866_out,
                 Y => SharedReg867_out);

   SharedReg868_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg867_out,
                 Y => SharedReg868_out);

   SharedReg869_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg868_out,
                 Y => SharedReg869_out);

   SharedReg870_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg869_out,
                 Y => SharedReg870_out);

   SharedReg871_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg870_out,
                 Y => SharedReg871_out);

   SharedReg872_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg871_out,
                 Y => SharedReg872_out);

   SharedReg873_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg872_out,
                 Y => SharedReg873_out);

   SharedReg874_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg873_out,
                 Y => SharedReg874_out);

   SharedReg875_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg874_out,
                 Y => SharedReg875_out);

   SharedReg876_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg875_out,
                 Y => SharedReg876_out);

   SharedReg877_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg876_out,
                 Y => SharedReg877_out);

   SharedReg878_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg877_out,
                 Y => SharedReg878_out);

   SharedReg879_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg878_out,
                 Y => SharedReg879_out);

   SharedReg880_instance: Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=28 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg879_out,
                 Y => SharedReg880_out);

   SharedReg881_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg880_out,
                 Y => SharedReg881_out);

   SharedReg882_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract3_6_impl_out,
                 Y => SharedReg882_out);

   SharedReg883_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg882_out,
                 Y => SharedReg883_out);

   SharedReg884_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg883_out,
                 Y => SharedReg884_out);

   SharedReg885_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg884_out,
                 Y => SharedReg885_out);

   SharedReg886_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg885_out,
                 Y => SharedReg886_out);

   SharedReg887_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg886_out,
                 Y => SharedReg887_out);

   SharedReg888_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg887_out,
                 Y => SharedReg888_out);

   SharedReg889_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg888_out,
                 Y => SharedReg889_out);

   SharedReg890_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg889_out,
                 Y => SharedReg890_out);

   SharedReg891_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg890_out,
                 Y => SharedReg891_out);

   SharedReg892_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg891_out,
                 Y => SharedReg892_out);

   SharedReg893_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg892_out,
                 Y => SharedReg893_out);

   SharedReg894_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg893_out,
                 Y => SharedReg894_out);

   SharedReg895_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg894_out,
                 Y => SharedReg895_out);

   SharedReg896_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg895_out,
                 Y => SharedReg896_out);

   SharedReg897_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg896_out,
                 Y => SharedReg897_out);

   SharedReg898_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg897_out,
                 Y => SharedReg898_out);

   SharedReg899_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg898_out,
                 Y => SharedReg899_out);

   SharedReg900_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg899_out,
                 Y => SharedReg900_out);

   SharedReg901_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg900_out,
                 Y => SharedReg901_out);

   SharedReg902_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg901_out,
                 Y => SharedReg902_out);

   SharedReg903_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg902_out,
                 Y => SharedReg903_out);

   SharedReg904_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg903_out,
                 Y => SharedReg904_out);

   SharedReg905_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg904_out,
                 Y => SharedReg905_out);

   SharedReg906_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract6_2_impl_out,
                 Y => SharedReg906_out);

   SharedReg907_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg906_out,
                 Y => SharedReg907_out);

   SharedReg908_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg907_out,
                 Y => SharedReg908_out);

   SharedReg909_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg908_out,
                 Y => SharedReg909_out);

   SharedReg910_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg909_out,
                 Y => SharedReg910_out);

   SharedReg911_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg910_out,
                 Y => SharedReg911_out);

   SharedReg912_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg911_out,
                 Y => SharedReg912_out);

   SharedReg913_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg912_out,
                 Y => SharedReg913_out);

   SharedReg914_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg913_out,
                 Y => SharedReg914_out);

   SharedReg915_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg914_out,
                 Y => SharedReg915_out);

   SharedReg916_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg915_out,
                 Y => SharedReg916_out);

   SharedReg917_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg916_out,
                 Y => SharedReg917_out);

   SharedReg918_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg917_out,
                 Y => SharedReg918_out);

   SharedReg919_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg918_out,
                 Y => SharedReg919_out);

   SharedReg920_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg919_out,
                 Y => SharedReg920_out);

   SharedReg921_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg920_out,
                 Y => SharedReg921_out);

   SharedReg922_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg921_out,
                 Y => SharedReg922_out);

   SharedReg923_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg922_out,
                 Y => SharedReg923_out);

   SharedReg924_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg923_out,
                 Y => SharedReg924_out);

   SharedReg925_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg924_out,
                 Y => SharedReg925_out);

   SharedReg926_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg925_out,
                 Y => SharedReg926_out);

   SharedReg927_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg926_out,
                 Y => SharedReg927_out);

   SharedReg928_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg927_out,
                 Y => SharedReg928_out);

   SharedReg929_instance: Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=28 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg928_out,
                 Y => SharedReg929_out);

   SharedReg930_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg929_out,
                 Y => SharedReg930_out);

   SharedReg931_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract6_4_impl_out,
                 Y => SharedReg931_out);

   SharedReg932_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg931_out,
                 Y => SharedReg932_out);

   SharedReg933_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg932_out,
                 Y => SharedReg933_out);

   SharedReg934_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg933_out,
                 Y => SharedReg934_out);

   SharedReg935_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg934_out,
                 Y => SharedReg935_out);

   SharedReg936_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg935_out,
                 Y => SharedReg936_out);

   SharedReg937_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg936_out,
                 Y => SharedReg937_out);

   SharedReg938_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg937_out,
                 Y => SharedReg938_out);

   SharedReg939_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg938_out,
                 Y => SharedReg939_out);

   SharedReg940_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg939_out,
                 Y => SharedReg940_out);

   SharedReg941_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg940_out,
                 Y => SharedReg941_out);

   SharedReg942_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg941_out,
                 Y => SharedReg942_out);

   SharedReg943_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg942_out,
                 Y => SharedReg943_out);

   SharedReg944_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg943_out,
                 Y => SharedReg944_out);

   SharedReg945_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg944_out,
                 Y => SharedReg945_out);

   SharedReg946_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg945_out,
                 Y => SharedReg946_out);

   SharedReg947_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg946_out,
                 Y => SharedReg947_out);

   SharedReg948_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg947_out,
                 Y => SharedReg948_out);

   SharedReg949_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg948_out,
                 Y => SharedReg949_out);

   SharedReg950_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg949_out,
                 Y => SharedReg950_out);

   SharedReg951_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg950_out,
                 Y => SharedReg951_out);

   SharedReg952_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg951_out,
                 Y => SharedReg952_out);

   SharedReg953_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg952_out,
                 Y => SharedReg953_out);

   SharedReg954_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg953_out,
                 Y => SharedReg954_out);

   SharedReg955_instance: Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=28 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg954_out,
                 Y => SharedReg955_out);

   SharedReg956_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg955_out,
                 Y => SharedReg956_out);

   SharedReg957_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract10_1_impl_out,
                 Y => SharedReg957_out);

   SharedReg958_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg957_out,
                 Y => SharedReg958_out);

   SharedReg959_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg958_out,
                 Y => SharedReg959_out);

   SharedReg960_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg959_out,
                 Y => SharedReg960_out);

   SharedReg961_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg960_out,
                 Y => SharedReg961_out);

   SharedReg962_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg961_out,
                 Y => SharedReg962_out);

   SharedReg963_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg962_out,
                 Y => SharedReg963_out);

   SharedReg964_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg963_out,
                 Y => SharedReg964_out);

   SharedReg965_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg964_out,
                 Y => SharedReg965_out);

   SharedReg966_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg965_out,
                 Y => SharedReg966_out);

   SharedReg967_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg966_out,
                 Y => SharedReg967_out);

   SharedReg968_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg967_out,
                 Y => SharedReg968_out);

   SharedReg969_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg968_out,
                 Y => SharedReg969_out);

   SharedReg970_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg969_out,
                 Y => SharedReg970_out);

   SharedReg971_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg970_out,
                 Y => SharedReg971_out);

   SharedReg972_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg971_out,
                 Y => SharedReg972_out);

   SharedReg973_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg972_out,
                 Y => SharedReg973_out);

   SharedReg974_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg973_out,
                 Y => SharedReg974_out);

   SharedReg975_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg974_out,
                 Y => SharedReg975_out);

   SharedReg976_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg975_out,
                 Y => SharedReg976_out);

   SharedReg977_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg976_out,
                 Y => SharedReg977_out);

   SharedReg978_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg977_out,
                 Y => SharedReg978_out);

   SharedReg979_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg978_out,
                 Y => SharedReg979_out);

   SharedReg980_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg979_out,
                 Y => SharedReg980_out);

   SharedReg981_instance: Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=28 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg980_out,
                 Y => SharedReg981_out);

   SharedReg982_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg981_out,
                 Y => SharedReg982_out);

   SharedReg983_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract12_6_impl_out,
                 Y => SharedReg983_out);

   SharedReg984_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg983_out,
                 Y => SharedReg984_out);

   SharedReg985_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg984_out,
                 Y => SharedReg985_out);

   SharedReg986_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg985_out,
                 Y => SharedReg986_out);

   SharedReg987_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg986_out,
                 Y => SharedReg987_out);

   SharedReg988_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg987_out,
                 Y => SharedReg988_out);

   SharedReg989_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg988_out,
                 Y => SharedReg989_out);

   SharedReg990_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg989_out,
                 Y => SharedReg990_out);

   SharedReg991_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg990_out,
                 Y => SharedReg991_out);

   SharedReg992_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg991_out,
                 Y => SharedReg992_out);

   SharedReg993_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg992_out,
                 Y => SharedReg993_out);

   SharedReg994_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg993_out,
                 Y => SharedReg994_out);

   SharedReg995_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg994_out,
                 Y => SharedReg995_out);

   SharedReg996_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg995_out,
                 Y => SharedReg996_out);

   SharedReg997_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg996_out,
                 Y => SharedReg997_out);

   SharedReg998_instance: Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=22 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg997_out,
                 Y => SharedReg998_out);

   SharedReg999_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg998_out,
                 Y => SharedReg999_out);

   SharedReg1000_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg999_out,
                 Y => SharedReg1000_out);

   SharedReg1001_instance: Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=28 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1000_out,
                 Y => SharedReg1001_out);

   SharedReg1002_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1001_out,
                 Y => SharedReg1002_out);

   SharedReg1003_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant2_0_impl_out,
                 Y => SharedReg1003_out);

   SharedReg1004_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1003_out,
                 Y => SharedReg1004_out);

   SharedReg1005_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1004_out,
                 Y => SharedReg1005_out);

   SharedReg1006_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1005_out,
                 Y => SharedReg1006_out);

   SharedReg1007_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1006_out,
                 Y => SharedReg1007_out);

   SharedReg1008_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1007_out,
                 Y => SharedReg1008_out);

   SharedReg1009_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1008_out,
                 Y => SharedReg1009_out);

   SharedReg1010_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1009_out,
                 Y => SharedReg1010_out);

   SharedReg1011_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1010_out,
                 Y => SharedReg1011_out);

   SharedReg1012_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1011_out,
                 Y => SharedReg1012_out);

   SharedReg1013_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1012_out,
                 Y => SharedReg1013_out);

   SharedReg1014_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1013_out,
                 Y => SharedReg1014_out);

   SharedReg1015_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1014_out,
                 Y => SharedReg1015_out);

   SharedReg1016_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1015_out,
                 Y => SharedReg1016_out);

   SharedReg1017_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1016_out,
                 Y => SharedReg1017_out);

   SharedReg1018_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1017_out,
                 Y => SharedReg1018_out);

   SharedReg1019_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1018_out,
                 Y => SharedReg1019_out);

   SharedReg1020_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1019_out,
                 Y => SharedReg1020_out);

   SharedReg1021_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1020_out,
                 Y => SharedReg1021_out);

   SharedReg1022_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1021_out,
                 Y => SharedReg1022_out);

   SharedReg1023_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1022_out,
                 Y => SharedReg1023_out);

   SharedReg1024_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1023_out,
                 Y => SharedReg1024_out);

   SharedReg1025_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1024_out,
                 Y => SharedReg1025_out);

   SharedReg1026_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1025_out,
                 Y => SharedReg1026_out);

   SharedReg1027_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1026_out,
                 Y => SharedReg1027_out);

   SharedReg1028_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1027_out,
                 Y => SharedReg1028_out);

   SharedReg1029_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1028_out,
                 Y => SharedReg1029_out);

   SharedReg1030_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1029_out,
                 Y => SharedReg1030_out);

   SharedReg1031_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1030_out,
                 Y => SharedReg1031_out);

   SharedReg1032_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1031_out,
                 Y => SharedReg1032_out);

   SharedReg1033_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1032_out,
                 Y => SharedReg1033_out);

   SharedReg1034_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1033_out,
                 Y => SharedReg1034_out);

   SharedReg1035_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1034_out,
                 Y => SharedReg1035_out);

   SharedReg1036_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1035_out,
                 Y => SharedReg1036_out);

   SharedReg1037_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1036_out,
                 Y => SharedReg1037_out);

   SharedReg1038_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1037_out,
                 Y => SharedReg1038_out);

   SharedReg1039_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1038_out,
                 Y => SharedReg1039_out);

   SharedReg1040_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1039_out,
                 Y => SharedReg1040_out);

   SharedReg1041_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1040_out,
                 Y => SharedReg1041_out);

   SharedReg1042_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1041_out,
                 Y => SharedReg1042_out);

   SharedReg1043_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1042_out,
                 Y => SharedReg1043_out);

   SharedReg1044_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1043_out,
                 Y => SharedReg1044_out);

   SharedReg1045_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1044_out,
                 Y => SharedReg1045_out);

   SharedReg1046_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1045_out,
                 Y => SharedReg1046_out);

   SharedReg1047_instance: Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=22 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1046_out,
                 Y => SharedReg1047_out);

   SharedReg1048_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1047_out,
                 Y => SharedReg1048_out);

   SharedReg1049_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1048_out,
                 Y => SharedReg1049_out);

   SharedReg1050_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1049_out,
                 Y => SharedReg1050_out);

   SharedReg1051_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1050_out,
                 Y => SharedReg1051_out);

   SharedReg1052_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1051_out,
                 Y => SharedReg1052_out);

   SharedReg1053_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1052_out,
                 Y => SharedReg1053_out);

   SharedReg1054_instance: Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=22 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1053_out,
                 Y => SharedReg1054_out);

   SharedReg1055_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1054_out,
                 Y => SharedReg1055_out);

   SharedReg1056_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1055_out,
                 Y => SharedReg1056_out);

   SharedReg1057_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant11_0_impl_out,
                 Y => SharedReg1057_out);

   SharedReg1058_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1057_out,
                 Y => SharedReg1058_out);

   SharedReg1059_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1058_out,
                 Y => SharedReg1059_out);

   SharedReg1060_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1059_out,
                 Y => SharedReg1060_out);

   SharedReg1061_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1060_out,
                 Y => SharedReg1061_out);

   SharedReg1062_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1061_out,
                 Y => SharedReg1062_out);

   SharedReg1063_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1062_out,
                 Y => SharedReg1063_out);

   SharedReg1064_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1063_out,
                 Y => SharedReg1064_out);

   SharedReg1065_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1064_out,
                 Y => SharedReg1065_out);

   SharedReg1066_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1065_out,
                 Y => SharedReg1066_out);

   SharedReg1067_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1066_out,
                 Y => SharedReg1067_out);

   SharedReg1068_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1067_out,
                 Y => SharedReg1068_out);

   SharedReg1069_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1068_out,
                 Y => SharedReg1069_out);

   SharedReg1070_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1069_out,
                 Y => SharedReg1070_out);

   SharedReg1071_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1070_out,
                 Y => SharedReg1071_out);

   SharedReg1072_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1071_out,
                 Y => SharedReg1072_out);

   SharedReg1073_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1072_out,
                 Y => SharedReg1073_out);

   SharedReg1074_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1073_out,
                 Y => SharedReg1074_out);

   SharedReg1075_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1074_out,
                 Y => SharedReg1075_out);

   SharedReg1076_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1075_out,
                 Y => SharedReg1076_out);

   SharedReg1077_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1076_out,
                 Y => SharedReg1077_out);

   SharedReg1078_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1077_out,
                 Y => SharedReg1078_out);

   SharedReg1079_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1078_out,
                 Y => SharedReg1079_out);

   SharedReg1080_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1079_out,
                 Y => SharedReg1080_out);

   SharedReg1081_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1080_out,
                 Y => SharedReg1081_out);

   SharedReg1082_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1081_out,
                 Y => SharedReg1082_out);

   SharedReg1083_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1082_out,
                 Y => SharedReg1083_out);

   SharedReg1084_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1083_out,
                 Y => SharedReg1084_out);

   SharedReg1085_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1084_out,
                 Y => SharedReg1085_out);

   SharedReg1086_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1085_out,
                 Y => SharedReg1086_out);

   SharedReg1087_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1086_out,
                 Y => SharedReg1087_out);

   SharedReg1088_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1087_out,
                 Y => SharedReg1088_out);

   SharedReg1089_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1088_out,
                 Y => SharedReg1089_out);

   SharedReg1090_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1089_out,
                 Y => SharedReg1090_out);

   SharedReg1091_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1090_out,
                 Y => SharedReg1091_out);

   SharedReg1092_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1091_out,
                 Y => SharedReg1092_out);

   SharedReg1093_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1092_out,
                 Y => SharedReg1093_out);

   SharedReg1094_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1093_out,
                 Y => SharedReg1094_out);

   SharedReg1095_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1094_out,
                 Y => SharedReg1095_out);

   SharedReg1096_instance: Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=22 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1095_out,
                 Y => SharedReg1096_out);

   SharedReg1097_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1096_out,
                 Y => SharedReg1097_out);

   SharedReg1098_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1097_out,
                 Y => SharedReg1098_out);

   SharedReg1099_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1098_out,
                 Y => SharedReg1099_out);

   SharedReg1100_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1099_out,
                 Y => SharedReg1100_out);

   SharedReg1101_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1100_out,
                 Y => SharedReg1101_out);

   SharedReg1102_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1101_out,
                 Y => SharedReg1102_out);

   SharedReg1103_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1102_out,
                 Y => SharedReg1103_out);

   SharedReg1104_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1103_out,
                 Y => SharedReg1104_out);

   SharedReg1105_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1104_out,
                 Y => SharedReg1105_out);

   SharedReg1106_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1105_out,
                 Y => SharedReg1106_out);

   SharedReg1107_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1106_out,
                 Y => SharedReg1107_out);

   SharedReg1108_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant4_0_impl_out,
                 Y => SharedReg1108_out);

   SharedReg1109_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1108_out,
                 Y => SharedReg1109_out);

   SharedReg1110_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1109_out,
                 Y => SharedReg1110_out);

   SharedReg1111_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1110_out,
                 Y => SharedReg1111_out);

   SharedReg1112_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1111_out,
                 Y => SharedReg1112_out);

   SharedReg1113_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1112_out,
                 Y => SharedReg1113_out);

   SharedReg1114_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant13_0_impl_out,
                 Y => SharedReg1114_out);

   SharedReg1115_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1114_out,
                 Y => SharedReg1115_out);

   SharedReg1116_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1115_out,
                 Y => SharedReg1116_out);

   SharedReg1117_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1116_out,
                 Y => SharedReg1117_out);

   SharedReg1118_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1117_out,
                 Y => SharedReg1118_out);

   SharedReg1119_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1118_out,
                 Y => SharedReg1119_out);

   SharedReg1120_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant5_0_impl_out,
                 Y => SharedReg1120_out);

   SharedReg1121_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant14_0_impl_out,
                 Y => SharedReg1121_out);

   SharedReg1122_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1121_out,
                 Y => SharedReg1122_out);

   SharedReg1123_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant6_0_impl_out,
                 Y => SharedReg1123_out);

   SharedReg1124_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1123_out,
                 Y => SharedReg1124_out);

   SharedReg1125_instance: Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=29 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1124_out,
                 Y => SharedReg1125_out);

   SharedReg1126_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1125_out,
                 Y => SharedReg1126_out);

   SharedReg1127_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1126_out,
                 Y => SharedReg1127_out);

   SharedReg1128_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1127_out,
                 Y => SharedReg1128_out);

   SharedReg1129_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1128_out,
                 Y => SharedReg1129_out);

   SharedReg1130_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1129_out,
                 Y => SharedReg1130_out);

   SharedReg1131_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1130_out,
                 Y => SharedReg1131_out);

   SharedReg1132_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1131_out,
                 Y => SharedReg1132_out);

   SharedReg1133_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1132_out,
                 Y => SharedReg1133_out);

   SharedReg1134_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1133_out,
                 Y => SharedReg1134_out);

   SharedReg1135_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1134_out,
                 Y => SharedReg1135_out);

   SharedReg1136_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant15_0_impl_out,
                 Y => SharedReg1136_out);

   SharedReg1137_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1136_out,
                 Y => SharedReg1137_out);

   SharedReg1138_instance: Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=29 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1137_out,
                 Y => SharedReg1138_out);

   SharedReg1139_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1138_out,
                 Y => SharedReg1139_out);

   SharedReg1140_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1139_out,
                 Y => SharedReg1140_out);

   SharedReg1141_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1140_out,
                 Y => SharedReg1141_out);

   SharedReg1142_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1141_out,
                 Y => SharedReg1142_out);

   SharedReg1143_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1142_out,
                 Y => SharedReg1143_out);

   SharedReg1144_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1143_out,
                 Y => SharedReg1144_out);

   SharedReg1145_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1144_out,
                 Y => SharedReg1145_out);

   SharedReg1146_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1145_out,
                 Y => SharedReg1146_out);

   SharedReg1147_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1146_out,
                 Y => SharedReg1147_out);

   SharedReg1148_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1147_out,
                 Y => SharedReg1148_out);

   SharedReg1149_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1148_out,
                 Y => SharedReg1149_out);

   SharedReg1150_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant7_0_impl_out,
                 Y => SharedReg1150_out);

   SharedReg1151_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1150_out,
                 Y => SharedReg1151_out);

   SharedReg1152_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant16_0_impl_out,
                 Y => SharedReg1152_out);

   SharedReg1153_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1152_out,
                 Y => SharedReg1153_out);

   SharedReg1154_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant8_0_impl_out,
                 Y => SharedReg1154_out);

   SharedReg1155_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1154_out,
                 Y => SharedReg1155_out);

   SharedReg1156_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1155_out,
                 Y => SharedReg1156_out);

   SharedReg1157_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1156_out,
                 Y => SharedReg1157_out);

   SharedReg1158_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1157_out,
                 Y => SharedReg1158_out);

   SharedReg1159_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1158_out,
                 Y => SharedReg1159_out);

   SharedReg1160_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant17_0_impl_out,
                 Y => SharedReg1160_out);

   SharedReg1161_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1160_out,
                 Y => SharedReg1161_out);

   SharedReg1162_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1161_out,
                 Y => SharedReg1162_out);

   SharedReg1163_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1162_out,
                 Y => SharedReg1163_out);

   SharedReg1164_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1163_out,
                 Y => SharedReg1164_out);

   SharedReg1165_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1164_out,
                 Y => SharedReg1165_out);

   SharedReg1166_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant9_0_impl_out,
                 Y => SharedReg1166_out);

   SharedReg1167_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1166_out,
                 Y => SharedReg1167_out);

   SharedReg1168_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant18_0_impl_out,
                 Y => SharedReg1168_out);

   SharedReg1169_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1168_out,
                 Y => SharedReg1169_out);

   SharedReg1170_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant_0_impl_out,
                 Y => SharedReg1170_out);

   SharedReg1171_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant1_0_impl_out,
                 Y => SharedReg1171_out);
end architecture;

