--------------------------------------------------------------------------------
--                         ModuloCounter_2_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity ModuloCounter_2_component is
   port ( clk, rst : in std_logic;
          Counter_out : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of ModuloCounter_2_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk,rst)
	 variable count : std_logic_vector(0 downto 0) := (others => '0');
begin
	 if rst = '1' then
	 	 count := (others => '0');
	 elsif clk'event and clk = '1' then
	 	 if count = 1 then
	 	 	 count := (others => '0');
	 	 else
	 	 	 count := count+1;
	 	 end if;
	 end if;
	 Counter_out <= count;
end process;
end architecture;

--------------------------------------------------------------------------------
--                          InputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2008)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity InputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(31 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of InputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal expInfty : std_logic := '0';
signal fracZero : std_logic := '0';
signal reprSubNormal : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal infinity : std_logic := '0';
signal zero : std_logic := '0';
signal NaN : std_logic := '0';
signal exnR : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   sX  <= X(31);
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   expInfty  <= '1' when expX = (7 downto 0 => '1') else '0';
   fracZero <= '1' when fracX = (22 downto 0 => '0') else '0';
   reprSubNormal <= fracX(22);
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= fracX(21 downto 0) & '0' when (expZero='1' and reprSubNormal='1')    else fracX;
   fracR <= sfracX;
   -- copy exponent. This will be OK even for subnormals, zero and infty since in such cases the exn bits will prevail
   expR <= expX;
   infinity <= expInfty and fracZero;
   zero <= expZero and not reprSubNormal;
   NaN <= expInfty and not fracZero;
   exnR <= 
           "00" when zero='1' 
      else "10" when infinity='1' 
      else "11" when NaN='1' 
      else "01" ;  -- normal number
   R <= exnR & sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--                         OutputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. Ferrandi  (2009-2012)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity OutputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of OutputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal exnX : std_logic_vector(1 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   exnX  <= X(33 downto 32);
   sX  <= X(31) when (exnX = "01" or exnX = "10" or exnX = "00") else '0';
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= 
      (22 downto 0 => '0') when (exnX = "00") else
      '1' & fracX(22 downto 1) when (expZero = '1' and exnX = "01") else
      fracX when (exnX = "01") else 
      (22 downto 1 => '0') & exnX(0);
   fracR <= sfracX;
   expR <=  
      (7 downto 0 => '0') when (exnX = "00") else
      expX when (exnX = "01") else 
      (7 downto 0 => '1');
   R <= sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      Y <= s0;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid391504_RightShifter
--                 (RightShifter_24_by_max_26_F250_uid391506)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid391504_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid391504_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_27_f250_uid391509
--                  (IntAdderAlternative_27_f250_uid391513)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid391509 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid391509 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--               LZCShifter_28_to_28_counting_32_F250_uid391516
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid391516 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid391516 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_34_f250_uid391519
--                   (IntAdderClassical_34_f250_uid391521)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid391519 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid391519 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                            FPAdd_8_23_uid391504
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid391504 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid391504 is
   component FPAdd_8_23_uid391504_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid391509 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid391516 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid391519 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid391504_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid391509  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid391516  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid391519  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   component FPAdd_8_23_uid391504 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= Y;
   FPAddSubOp_instance: FPAdd_8_23_uid391504  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_2_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_2_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(0 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_2_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "0",
         iS_1 when "1",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--          IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid392594
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid392594 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          Y : in std_logic_vector(23 downto 0);
          R : out std_logic_vector(47 downto 0)   );
end entity;

architecture arch of IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid392594 is
signal XX_m392595 : std_logic_vector(23 downto 0) := (others => '0');
signal YY_m392595 : std_logic_vector(23 downto 0) := (others => '0');
signal XX : unsigned(-1+24 downto 0) := (others => '0');
signal YY : unsigned(-1+24 downto 0) := (others => '0');
signal RR : unsigned(-1+48 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   XX_m392595 <= X ;
   YY_m392595 <= Y ;
   XX <= unsigned(X);
   YY <= unsigned(Y);
   RR <= XX*YY;
   R <= std_logic_vector(RR(47 downto 0));
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_33_f500_uid392598
--                   (IntAdderClassical_33_f500_uid392600)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_33_f500_uid392598 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(32 downto 0);
          Y : in std_logic_vector(32 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(32 downto 0)   );
end entity;

architecture arch of IntAdder_33_f500_uid392598 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--         FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin 2008-2011
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   component IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid392594 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             Y : in std_logic_vector(23 downto 0);
             R : out std_logic_vector(47 downto 0)   );
   end component;

   component IntAdder_33_f500_uid392598 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(32 downto 0);
             Y : in std_logic_vector(32 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(32 downto 0)   );
   end component;

signal sign, sign_d1, sign_d2 : std_logic := '0';
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal expY : std_logic_vector(7 downto 0) := (others => '0');
signal expSumPreSub, expSumPreSub_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal bias, bias_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal expSum : std_logic_vector(9 downto 0) := (others => '0');
signal sigX : std_logic_vector(23 downto 0) := (others => '0');
signal sigY : std_logic_vector(23 downto 0) := (others => '0');
signal sigProd, sigProd_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal excSel : std_logic_vector(3 downto 0) := (others => '0');
signal exc, exc_d1, exc_d2 : std_logic_vector(1 downto 0) := (others => '0');
signal norm : std_logic := '0';
signal expPostNorm : std_logic_vector(9 downto 0) := (others => '0');
signal sigProdExt, sigProdExt_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal expSig, expSig_d1 : std_logic_vector(32 downto 0) := (others => '0');
signal sticky, sticky_d1 : std_logic := '0';
signal guard, guard_d1 : std_logic := '0';
signal round : std_logic := '0';
signal expSigPostRound : std_logic_vector(32 downto 0) := (others => '0');
signal excPostNorm : std_logic_vector(1 downto 0) := (others => '0');
signal finalExc : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            sign_d1 <=  sign;
            sign_d2 <=  sign_d1;
            expSumPreSub_d1 <=  expSumPreSub;
            bias_d1 <=  bias;
            sigProd_d1 <=  sigProd;
            exc_d1 <=  exc;
            exc_d2 <=  exc_d1;
            sigProdExt_d1 <=  sigProdExt;
            expSig_d1 <=  expSig;
            sticky_d1 <=  sticky;
            guard_d1 <=  guard;
         end if;
      end process;
   sign <= X(31) xor Y(31);
   expX <= X(30 downto 23);
   expY <= Y(30 downto 23);
   expSumPreSub <= ("00" & expX) + ("00" & expY);
   bias <= CONV_STD_LOGIC_VECTOR(127,10);
   ----------------Synchro barrier, entering cycle 1----------------
   expSum <= expSumPreSub_d1 - bias_d1;
   ----------------Synchro barrier, entering cycle 0----------------
   sigX <= "1" & X(22 downto 0);
   sigY <= "1" & Y(22 downto 0);
   SignificandMultiplication: IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid392594  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => sigProd,
                 X => sigX,
                 Y => sigY);
   ----------------Synchro barrier, entering cycle 0----------------
   excSel <= X(33 downto 32) & Y(33 downto 32);
   with excSel select 
   exc <= "00" when  "0000" | "0001" | "0100", 
          "01" when "0101",
          "10" when "0110" | "1001" | "1010" ,
          "11" when others;
   norm <= sigProd_d1(47);
   -- exponent update
   expPostNorm <= expSum + ("000000000" & norm);
   -- significand normalization shift
   sigProdExt <= sigProd_d1(46 downto 0) & "0" when norm='1' else
                         sigProd_d1(45 downto 0) & "00";
   expSig <= expPostNorm & sigProdExt(47 downto 25);
   sticky <= sigProdExt(24);
   guard <= '0' when sigProdExt(23 downto 0)="000000000000000000000000" else '1';
   ----------------Synchro barrier, entering cycle 2----------------
   round <= sticky_d1 and ( (guard_d1 and not(sigProdExt_d1(25))) or (sigProdExt_d1(25) ))  ;
   RoundingAdder: IntAdder_33_f500_uid392598  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => round,
                 R => expSigPostRound   ,
                 X => expSig_d1,
                 Y => "000000000000000000000000000000000");
   with expSigPostRound(32 downto 31) select
   excPostNorm <=  "01"  when  "00",
                               "10"             when "01", 
                               "00"             when "11"|"10",
                               "11"             when others;
   with exc_d2 select 
   finalExc <= exc_d2 when  "11"|"10"|"00",
                       excPostNorm when others; 
   R <= finalExc & sign_d2 & expSigPostRound(30 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid392681_RightShifter
--                 (RightShifter_24_by_max_26_F250_uid392683)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid392681_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid392681_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_27_f250_uid392686
--                  (IntAdderAlternative_27_f250_uid392690)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid392686 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid392686 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--               LZCShifter_28_to_28_counting_32_F250_uid392693
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid392693 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid392693 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_34_f250_uid392696
--                   (IntAdderClassical_34_f250_uid392698)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid392696 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid392696 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                            FPAdd_8_23_uid392681
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid392681 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid392681 is
   component FPAdd_8_23_uid392681_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid392686 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid392693 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid392696 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid392681_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid392686  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid392693  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid392696  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
   component FPAdd_8_23_uid392681 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= (Y(Y'length-1 downto Y'length-2)) & (not Y(Y'length-3)) & Y(Y'length-4 downto 0);
   FPAddSubOp_instance: FPAdd_8_23_uid392681  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--                      Constant_float_8_23_1_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_1_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_1_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111100000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                      Constant_float_8_23_0_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_0_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_0_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0000000000000000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_cosnpi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosnpi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosnpi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_sinnpi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinnpi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinnpi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn3_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn3_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn3_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn3_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn3_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn3_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_cosnpi_div_2_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosnpi_div_2_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosnpi_div_2_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0000000000000000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_sinnpi_div_2_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinnpi_div_2_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinnpi_div_2_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111100000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn5_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn5_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn5_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn5_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn5_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn5_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn3_mult_pi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn3_mult_pi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn3_mult_pi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn3_mult_pi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn3_mult_pi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn3_mult_pi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn7_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn7_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn7_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn7_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn7_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn7_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_cosnpi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosnpi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosnpi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_sinnpi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinnpi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinnpi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 7 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      Y <= s6;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      Y <= s5;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 20 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      Y <= s19;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 21 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      Y <= s20;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 35 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      Y <= s34;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                         implementedSystem_toplevel
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity implementedSystem_toplevel is
   port ( clk, rst : in std_logic;
          x0_re : in std_logic_vector(31 downto 0);
          x0_im : in std_logic_vector(31 downto 0);
          x1_re : in std_logic_vector(31 downto 0);
          x1_im : in std_logic_vector(31 downto 0);
          x2_re : in std_logic_vector(31 downto 0);
          x2_im : in std_logic_vector(31 downto 0);
          x3_re : in std_logic_vector(31 downto 0);
          x3_im : in std_logic_vector(31 downto 0);
          x4_re : in std_logic_vector(31 downto 0);
          x4_im : in std_logic_vector(31 downto 0);
          x5_re : in std_logic_vector(31 downto 0);
          x5_im : in std_logic_vector(31 downto 0);
          x6_re : in std_logic_vector(31 downto 0);
          x6_im : in std_logic_vector(31 downto 0);
          x7_re : in std_logic_vector(31 downto 0);
          x7_im : in std_logic_vector(31 downto 0);
          x8_re : in std_logic_vector(31 downto 0);
          x8_im : in std_logic_vector(31 downto 0);
          x9_re : in std_logic_vector(31 downto 0);
          x9_im : in std_logic_vector(31 downto 0);
          x10_re : in std_logic_vector(31 downto 0);
          x10_im : in std_logic_vector(31 downto 0);
          x11_re : in std_logic_vector(31 downto 0);
          x11_im : in std_logic_vector(31 downto 0);
          x12_re : in std_logic_vector(31 downto 0);
          x12_im : in std_logic_vector(31 downto 0);
          x13_re : in std_logic_vector(31 downto 0);
          x13_im : in std_logic_vector(31 downto 0);
          x14_re : in std_logic_vector(31 downto 0);
          x14_im : in std_logic_vector(31 downto 0);
          x15_re : in std_logic_vector(31 downto 0);
          x15_im : in std_logic_vector(31 downto 0);
          y0_re : out std_logic_vector(31 downto 0);
          y0_im : out std_logic_vector(31 downto 0);
          y1_re : out std_logic_vector(31 downto 0);
          y1_im : out std_logic_vector(31 downto 0);
          y2_re : out std_logic_vector(31 downto 0);
          y2_im : out std_logic_vector(31 downto 0);
          y3_re : out std_logic_vector(31 downto 0);
          y3_im : out std_logic_vector(31 downto 0);
          y4_re : out std_logic_vector(31 downto 0);
          y4_im : out std_logic_vector(31 downto 0);
          y5_re : out std_logic_vector(31 downto 0);
          y5_im : out std_logic_vector(31 downto 0);
          y6_re : out std_logic_vector(31 downto 0);
          y6_im : out std_logic_vector(31 downto 0);
          y7_re : out std_logic_vector(31 downto 0);
          y7_im : out std_logic_vector(31 downto 0);
          y8_re : out std_logic_vector(31 downto 0);
          y8_im : out std_logic_vector(31 downto 0);
          y9_re : out std_logic_vector(31 downto 0);
          y9_im : out std_logic_vector(31 downto 0);
          y10_re : out std_logic_vector(31 downto 0);
          y10_im : out std_logic_vector(31 downto 0);
          y11_re : out std_logic_vector(31 downto 0);
          y11_im : out std_logic_vector(31 downto 0);
          y12_re : out std_logic_vector(31 downto 0);
          y12_im : out std_logic_vector(31 downto 0);
          y13_re : out std_logic_vector(31 downto 0);
          y13_im : out std_logic_vector(31 downto 0);
          y14_re : out std_logic_vector(31 downto 0);
          y14_im : out std_logic_vector(31 downto 0);
          y15_re : out std_logic_vector(31 downto 0);
          y15_im : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of implementedSystem_toplevel is
   component ModuloCounter_2_component is
      port ( clk, rst : in std_logic;
             Counter_out : out std_logic_vector(0 downto 0)   );
   end component;

   component InputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(31 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component OutputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(31 downto 0)   );
   end component;

   component Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_2_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(0 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_1_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_0_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosnpi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinnpi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn3_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn3_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosnpi_div_2_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinnpi_div_2_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn5_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn5_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn3_mult_pi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn3_mult_pi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn7_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn7_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosnpi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinnpi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

signal ModCount21_out : std_logic_vector(0 downto 0) := (others => '0');
signal x0_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x0_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x1_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x1_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x2_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x2_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x3_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x3_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x4_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x4_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x5_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x5_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x6_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x6_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x7_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x7_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x8_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x8_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x9_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x9_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x10_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x10_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x11_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x11_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x12_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x12_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x13_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x13_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x14_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x14_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x15_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x15_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No14_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No15_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No16_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No17_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No18_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No19_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No20_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No21_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No22_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No23_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No24_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No25_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No26_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No27_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No28_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No29_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No30_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No31_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No32_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No33_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No34_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No35_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add12_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No36_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No37_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add13_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add13_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No38_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add13_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No39_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add14_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add14_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No40_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add14_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No41_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No42_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No43_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add15_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add15_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No44_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add15_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No45_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add7_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add7_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No46_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add7_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No47_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add16_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add16_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No48_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add16_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No49_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add8_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add8_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No50_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add8_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No51_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add9_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add9_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No52_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add9_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No53_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add18_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add18_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No54_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add18_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No55_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add20_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add20_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No56_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add20_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No57_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add110_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add110_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No58_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add110_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No59_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add22_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add22_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No60_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add22_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No61_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add112_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add112_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No62_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add112_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No63_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add24_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add24_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No64_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add24_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No65_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add114_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add114_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No66_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add114_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No67_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add25_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add25_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No68_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add25_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No69_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add115_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add115_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No70_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add115_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No71_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add26_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add26_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No72_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add26_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No73_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add116_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add116_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No74_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add116_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No75_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add27_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add27_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No76_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add27_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No77_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add117_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add117_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No78_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add117_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No79_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add34_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add34_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No80_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add34_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No81_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add124_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add124_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No82_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add124_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No83_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add126_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add126_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No84_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add126_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No85_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add37_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add37_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No86_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add37_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No87_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add127_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add127_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No88_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add127_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No89_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add129_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add129_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No90_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add129_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No91_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add41_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add41_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No92_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add41_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No93_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add131_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add131_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No94_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add131_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No95_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add43_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add43_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No96_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add43_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No97_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No98_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No99_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product11_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No100_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No101_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No102_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No103_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product31_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No104_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No105_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No106_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No107_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No108_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No109_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No110_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No111_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add45_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add45_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No112_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add45_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No113_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No114_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No115_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product13_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product13_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No116_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product13_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No117_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product23_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No118_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No119_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product33_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No120_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No121_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No122_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No123_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add46_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add46_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No124_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add46_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No125_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product7_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product7_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No126_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product7_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No127_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product14_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product14_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No128_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product14_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No129_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product24_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product24_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No130_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product24_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No131_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add47_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add47_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No132_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add47_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No133_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product8_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product8_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No134_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product8_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No135_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product15_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product15_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No136_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product15_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No137_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product25_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product25_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No138_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product25_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No139_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product35_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product35_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No140_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product35_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No141_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No142_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No143_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add48_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add48_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No144_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add48_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No145_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product9_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product9_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No146_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product9_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No147_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product16_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product16_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No148_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product16_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No149_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product26_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product26_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No150_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product26_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No151_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product36_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product36_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No152_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product36_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No153_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract7_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract7_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No154_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract7_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No155_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add49_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add49_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No156_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add49_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No157_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product10_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product10_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No158_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product10_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No159_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product17_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product17_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No160_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product17_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No161_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product27_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product27_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No162_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product27_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No163_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product37_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product37_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No164_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product37_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No165_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract8_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract8_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No166_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract8_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No167_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add50_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add50_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No168_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add50_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No169_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product18_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product18_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No170_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product18_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No171_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product19_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product19_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No172_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product19_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No173_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product28_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No174_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No175_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product38_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product38_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No176_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product38_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No177_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract9_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No178_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No179_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add52_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add52_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No180_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add52_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No181_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product30_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product30_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No182_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product30_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No183_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product111_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No184_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No185_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product210_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No186_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No187_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product310_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No188_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No189_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract11_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract11_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No190_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract11_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No191_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add53_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add53_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No192_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add53_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No193_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product40_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product40_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No194_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product40_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No195_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product112_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product112_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No196_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product112_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No197_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product211_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product211_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No198_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product211_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No199_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product311_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product311_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No200_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product311_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No201_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract12_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No202_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No203_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add54_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add54_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No204_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add54_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No205_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product41_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product41_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No206_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product41_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No207_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product113_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product113_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No208_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product113_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No209_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product212_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product212_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No210_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product212_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No211_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product312_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product312_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No212_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product312_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No213_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract13_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract13_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No214_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract13_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No215_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add56_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add56_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No216_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add56_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No217_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product43_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product43_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No218_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product43_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No219_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product115_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product115_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No220_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product115_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No221_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product214_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product214_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No222_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product214_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No223_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product314_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product314_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No224_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product314_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No225_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract15_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract15_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No226_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract15_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No227_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add57_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add57_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No228_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add57_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No229_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product44_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product44_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No230_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product44_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No231_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product116_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product116_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No232_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product116_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No233_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product215_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product215_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No234_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product215_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No235_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product315_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product315_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No236_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product315_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No237_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract16_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract16_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No238_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract16_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No239_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add58_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add58_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No240_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add58_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No241_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product45_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product45_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No242_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product45_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No243_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product117_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product117_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No244_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product117_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No245_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product216_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product216_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No246_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product216_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No247_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product316_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product316_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No248_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product316_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No249_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract17_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract17_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No250_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract17_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No251_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add59_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add59_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No252_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add59_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No253_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product46_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product46_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No254_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product46_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No255_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product118_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product118_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No256_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product118_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No257_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product217_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product217_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No258_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product217_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No259_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product317_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product317_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No260_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product317_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No261_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract18_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract18_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No262_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract18_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No263_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add61_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add61_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No264_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add61_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No265_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product48_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product48_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No266_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product48_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No267_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product120_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product120_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No268_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product120_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No269_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product219_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product219_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No270_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product219_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No271_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product319_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product319_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No272_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product319_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No273_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract20_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract20_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No274_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract20_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No275_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add63_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add63_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No276_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add63_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No277_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product50_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product50_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No278_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product50_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No279_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product122_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product122_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No280_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product122_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No281_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product221_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product221_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No282_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product221_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No283_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product321_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No284_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No285_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract22_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract22_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No286_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract22_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No287_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add65_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add65_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No288_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add65_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No289_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product52_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product52_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No290_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product52_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No291_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product124_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product124_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No292_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product124_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No293_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product223_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product223_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No294_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product223_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No295_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product323_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product323_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No296_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product323_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No297_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract24_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract24_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No298_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract24_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No299_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add66_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add66_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No300_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add66_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No301_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product53_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product53_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No302_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product53_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No303_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product125_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product125_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No304_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product125_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No305_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product224_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product224_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No306_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product224_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No307_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product324_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product324_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No308_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product324_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No309_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract25_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract25_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No310_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract25_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No311_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add67_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add67_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No312_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add67_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No313_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product54_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product54_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No314_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product54_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No315_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product126_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product126_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No316_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product126_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No317_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product225_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product225_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No318_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product225_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No319_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product325_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product325_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No320_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product325_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No321_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract26_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract26_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No322_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract26_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No323_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add68_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add68_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No324_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add68_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No325_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product55_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product55_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No326_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product55_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No327_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product127_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product127_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No328_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product127_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No329_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product226_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product226_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No330_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product226_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No331_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product326_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product326_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No332_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product326_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No333_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract27_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract27_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No334_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract27_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No335_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add83_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add83_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No336_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add83_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No337_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product70_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product70_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No338_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product70_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No339_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product142_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product142_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No340_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product142_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No341_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product241_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product241_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No342_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product241_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No343_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product341_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product341_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No344_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product341_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No345_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract42_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract42_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No346_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract42_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No347_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add84_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add84_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No348_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add84_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No349_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product71_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product71_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No350_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product71_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No351_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product143_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product143_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No352_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product143_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No353_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product242_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product242_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No354_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product242_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No355_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product342_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product342_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No356_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product342_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No357_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract43_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract43_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No358_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract43_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No359_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add85_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add85_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No360_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add85_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No361_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product72_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product72_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No362_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product72_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No363_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product144_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product144_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No364_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product144_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No365_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product243_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product243_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No366_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product243_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No367_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product343_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product343_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No368_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product343_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No369_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract44_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract44_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No370_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract44_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No371_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract45_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract45_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No372_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract45_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No373_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add87_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add87_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No374_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add87_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No375_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product74_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product74_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No376_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product74_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No377_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product146_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product146_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No378_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product146_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No379_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product245_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product245_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No380_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product245_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No381_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product345_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product345_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No382_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product345_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No383_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract46_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract46_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No384_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract46_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No385_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract47_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract47_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No386_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract47_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No387_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract48_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract48_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No388_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract48_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No389_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract49_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract49_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No390_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract49_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No391_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract50_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract50_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No392_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract50_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No393_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract52_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract52_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No394_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract52_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No395_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract112_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract112_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No396_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract112_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No397_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract114_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract114_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No398_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract114_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No399_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract55_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract55_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No400_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract55_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No401_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract115_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract115_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No402_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract115_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No403_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract56_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract56_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No404_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract56_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No405_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract116_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract116_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No406_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract116_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No407_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract57_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract57_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No408_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract57_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No409_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract117_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract117_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No410_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract117_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No411_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract59_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract59_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No412_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract59_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No413_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract119_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract119_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No414_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract119_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No415_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract62_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract62_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No416_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract62_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No417_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract122_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract122_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No418_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract122_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No419_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract63_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract63_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No420_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract63_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No421_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract123_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract123_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No422_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract123_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No423_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract127_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract127_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No424_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract127_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No425_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract68_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract68_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No426_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract68_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No427_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract71_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract71_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No428_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract71_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No429_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract131_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract131_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No430_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract131_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No431_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract72_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract72_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No432_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract72_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No433_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract132_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract132_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No434_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract132_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No435_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract74_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract74_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No436_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract74_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No437_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract134_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract134_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No438_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract134_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No439_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract75_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract75_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No440_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract75_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No441_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract135_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract135_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No442_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract135_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No443_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract80_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract80_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No444_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract80_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No445_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract140_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract140_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No446_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract140_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No447_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant11_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant12_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant13_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant14_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant15_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant7_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant16_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant8_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant17_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant9_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant18_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant10_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant19_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant20_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant110_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant21_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant111_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant22_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant112_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant23_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant113_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant24_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant114_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant25_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant115_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant26_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant116_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant27_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant117_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant28_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant118_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant29_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant119_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant30_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant120_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant31_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant121_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant32_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant122_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant33_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant123_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant34_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant124_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant35_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant125_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant36_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant126_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant37_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant127_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant38_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant128_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant39_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant129_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant40_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant130_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant41_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant131_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant42_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant132_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant43_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant133_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant44_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant134_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant45_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant135_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant46_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant136_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant47_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant137_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant48_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant138_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant49_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant139_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant50_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant140_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant51_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant141_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant52_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant142_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant53_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant143_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant54_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant144_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant55_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant145_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant56_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant146_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant57_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant147_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No14_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No15_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No40_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No41_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No42_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No43_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No44_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No45_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No46_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No47_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No48_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No49_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No50_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No51_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No52_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No53_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No54_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No55_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out : std_logic_vector(33 downto 0) := (others => '0');
signal x0_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x0_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x1_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x1_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x2_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x2_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x3_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x3_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x4_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x4_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x5_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x5_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x6_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x6_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x7_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x7_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x8_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x8_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x9_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x9_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x10_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x10_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x11_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x11_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x12_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x12_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x13_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x13_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x14_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x14_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x15_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x15_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y0_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y0_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y1_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y1_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y2_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y2_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y3_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y3_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y4_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y4_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y5_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y5_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y6_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y6_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y7_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y7_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y8_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y8_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y9_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y9_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y10_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y10_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y11_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y11_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y12_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y12_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y13_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y13_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y14_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y14_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y15_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y15_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Delay1No32_out_to_Add2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No33_out_to_Add2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No8_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No34_out_to_Add11_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No35_out_to_Add11_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No1_out_to_MUX_Add11_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add11_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No9_out_to_MUX_Add11_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add11_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No36_out_to_Add12_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No37_out_to_Add12_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Add12_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add12_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Add12_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add12_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No38_out_to_Add13_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No39_out_to_Add13_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Add13_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Add13_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Add13_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Add13_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No40_out_to_Add14_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No41_out_to_Add14_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Add14_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Add14_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Add14_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Add14_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No42_out_to_Add6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No43_out_to_Add6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Add6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Add6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Add6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Add6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No44_out_to_Add15_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No45_out_to_Add15_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Add15_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Add15_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Add15_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Add15_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No46_out_to_Add7_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No47_out_to_Add7_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No48_out_to_Add16_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No49_out_to_Add16_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No2_out_to_MUX_Add16_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Add16_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No10_out_to_MUX_Add16_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Add16_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No50_out_to_Add8_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No51_out_to_Add8_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No3_out_to_MUX_Add8_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Add8_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No11_out_to_MUX_Add8_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Add8_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No52_out_to_Add9_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No53_out_to_Add9_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No54_out_to_Add18_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No55_out_to_Add18_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Add18_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Add18_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Add18_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Add18_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No56_out_to_Add20_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No57_out_to_Add20_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Add20_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Add20_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Add20_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Add20_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No58_out_to_Add110_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No59_out_to_Add110_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Add110_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Add110_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Add110_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Add110_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No60_out_to_Add22_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No61_out_to_Add22_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Add22_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Add22_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Add22_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Add22_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No62_out_to_Add112_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No63_out_to_Add112_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Add112_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Add112_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Add112_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Add112_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No64_out_to_Add24_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No65_out_to_Add24_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Add24_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Add24_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Add24_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Add24_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No66_out_to_Add114_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No67_out_to_Add114_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Add114_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Add114_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Add114_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Add114_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No68_out_to_Add25_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No69_out_to_Add25_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Add25_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Add25_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Add25_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Add25_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No70_out_to_Add115_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No71_out_to_Add115_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Add115_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Add115_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Add115_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Add115_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No72_out_to_Add26_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No73_out_to_Add26_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Add26_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Add26_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Add26_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Add26_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No74_out_to_Add116_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No75_out_to_Add116_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Add116_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Add116_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Add116_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Add116_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No76_out_to_Add27_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No77_out_to_Add27_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No6_out_to_MUX_Add27_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Add27_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No14_out_to_MUX_Add27_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Add27_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No78_out_to_Add117_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No79_out_to_Add117_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Add117_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Add117_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out_to_MUX_Add117_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Add117_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No80_out_to_Add34_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No81_out_to_Add34_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Add34_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Add34_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out_to_MUX_Add34_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add34_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No82_out_to_Add124_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No83_out_to_Add124_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out_to_MUX_Add124_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add124_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Add124_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add124_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No84_out_to_Add126_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No85_out_to_Add126_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Add126_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add126_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Add126_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add126_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No86_out_to_Add37_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No87_out_to_Add37_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No4_out_to_MUX_Add37_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add37_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No12_out_to_MUX_Add37_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add37_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No88_out_to_Add127_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No89_out_to_Add127_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No5_out_to_MUX_Add127_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Add127_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No13_out_to_MUX_Add127_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add127_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No90_out_to_Add129_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No91_out_to_Add129_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No7_out_to_MUX_Add129_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add129_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No15_out_to_MUX_Add129_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add129_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No92_out_to_Add41_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No93_out_to_Add41_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Add41_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Add41_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Add41_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Add41_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No94_out_to_Add131_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No95_out_to_Add131_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Add131_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Add131_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Add131_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out_to_MUX_Add131_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No96_out_to_Add43_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No97_out_to_Add43_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_Add43_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Add43_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Add43_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_Add43_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No98_out_to_Product4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No99_out_to_Product4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No100_out_to_Product11_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No101_out_to_Product11_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Product11_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Product11_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product11_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product11_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No102_out_to_Product21_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No103_out_to_Product21_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No104_out_to_Product31_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No105_out_to_Product31_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Product31_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product31_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product31_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Product31_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No106_out_to_Subtract2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No107_out_to_Subtract2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No108_out_to_Product32_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No109_out_to_Product32_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product32_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Product32_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Product32_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product32_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No110_out_to_Subtract3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No111_out_to_Subtract3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Subtract3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Subtract3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Subtract3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Subtract3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No112_out_to_Add45_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No113_out_to_Add45_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Add45_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Add45_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Add45_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Add45_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No114_out_to_Product6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No115_out_to_Product6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Product6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Product6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Product6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No116_out_to_Product13_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No117_out_to_Product13_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No118_out_to_Product23_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No119_out_to_Product23_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No120_out_to_Product33_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No121_out_to_Product33_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No122_out_to_Subtract4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No123_out_to_Subtract4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No124_out_to_Add46_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No125_out_to_Add46_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Add46_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Add46_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Add46_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Add46_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No126_out_to_Product7_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No127_out_to_Product7_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No128_out_to_Product14_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No129_out_to_Product14_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Product14_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Product14_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Product14_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product14_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No130_out_to_Product24_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No131_out_to_Product24_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Product24_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Product24_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Product24_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product24_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No132_out_to_Add47_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No133_out_to_Add47_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Add47_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Add47_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Add47_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Add47_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No134_out_to_Product8_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No135_out_to_Product8_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Product8_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Product8_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Product8_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product8_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No136_out_to_Product15_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No137_out_to_Product15_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Product15_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product15_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Product15_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Product15_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No138_out_to_Product25_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No139_out_to_Product25_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Product25_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Product25_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Product25_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product25_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No140_out_to_Product35_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No141_out_to_Product35_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Product35_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Product35_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Product35_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product35_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No142_out_to_Subtract6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No143_out_to_Subtract6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Subtract6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Subtract6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Subtract6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Subtract6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No144_out_to_Add48_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No145_out_to_Add48_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Add48_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Add48_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Add48_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Add48_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No146_out_to_Product9_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No147_out_to_Product9_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Product9_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Product9_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Product9_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out_to_MUX_Product9_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No148_out_to_Product16_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No149_out_to_Product16_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Product16_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Product16_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Product16_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Product16_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No150_out_to_Product26_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No151_out_to_Product26_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Product26_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Product26_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Product26_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out_to_MUX_Product26_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No152_out_to_Product36_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No153_out_to_Product36_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Product36_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Product36_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Product36_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Product36_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No154_out_to_Subtract7_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No155_out_to_Subtract7_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Subtract7_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Subtract7_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Subtract7_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Subtract7_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No156_out_to_Add49_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No157_out_to_Add49_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Add49_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Add49_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Add49_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Add49_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No158_out_to_Product10_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No159_out_to_Product10_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Product10_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Product10_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Product10_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Product10_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No160_out_to_Product17_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No161_out_to_Product17_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Product17_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Product17_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Product17_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Product17_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No162_out_to_Product27_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No163_out_to_Product27_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Product27_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Product27_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Product27_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Product27_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No164_out_to_Product37_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No165_out_to_Product37_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Product37_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out_to_MUX_Product37_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Product37_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Product37_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No166_out_to_Subtract8_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No167_out_to_Subtract8_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Subtract8_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Subtract8_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Subtract8_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Subtract8_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No168_out_to_Add50_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No169_out_to_Add50_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Add50_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Add50_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Add50_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Add50_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No170_out_to_Product18_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No171_out_to_Product18_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out_to_MUX_Product18_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out_to_MUX_Product18_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Product18_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out_to_MUX_Product18_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No172_out_to_Product19_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No173_out_to_Product19_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out_to_MUX_Product19_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Product19_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out_to_MUX_Product19_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Product19_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No174_out_to_Product28_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No175_out_to_Product28_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Product28_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out_to_MUX_Product28_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Product28_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Product28_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No176_out_to_Product38_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No177_out_to_Product38_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out_to_MUX_Product38_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Product38_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Product38_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product38_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No178_out_to_Subtract9_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No179_out_to_Subtract9_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Subtract9_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Subtract9_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Subtract9_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Subtract9_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No180_out_to_Add52_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No181_out_to_Add52_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Add52_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Add52_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Add52_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Add52_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No182_out_to_Product30_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No183_out_to_Product30_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Product30_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Product30_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product30_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product30_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No184_out_to_Product111_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No185_out_to_Product111_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Product111_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Product111_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product111_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product111_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No186_out_to_Product210_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No187_out_to_Product210_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Product210_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product210_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product210_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Product210_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No188_out_to_Product310_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No189_out_to_Product310_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product310_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out_to_MUX_Product310_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Product310_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Product310_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No190_out_to_Subtract11_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No191_out_to_Subtract11_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Subtract11_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Subtract11_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Subtract11_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Subtract11_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No192_out_to_Add53_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No193_out_to_Add53_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Add53_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Add53_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Add53_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Add53_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No194_out_to_Product40_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No195_out_to_Product40_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Product40_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out_to_MUX_Product40_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product40_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Product40_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No196_out_to_Product112_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No197_out_to_Product112_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Product112_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Product112_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product112_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Product112_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No198_out_to_Product211_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No199_out_to_Product211_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Product211_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Product211_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product211_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Product211_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No200_out_to_Product311_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No201_out_to_Product311_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product311_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Product311_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Product311_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Product311_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No202_out_to_Subtract12_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No203_out_to_Subtract12_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Subtract12_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Subtract12_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Subtract12_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Subtract12_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No204_out_to_Add54_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No205_out_to_Add54_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Add54_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Add54_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Add54_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Add54_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No206_out_to_Product41_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No207_out_to_Product41_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out_to_MUX_Product41_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Product41_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product41_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product41_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No208_out_to_Product113_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No209_out_to_Product113_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out_to_MUX_Product113_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Product113_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product113_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product113_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No210_out_to_Product212_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No211_out_to_Product212_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out_to_MUX_Product212_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Product212_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product212_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product212_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No212_out_to_Product312_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No213_out_to_Product312_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product312_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product312_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out_to_MUX_Product312_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Product312_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No214_out_to_Subtract13_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No215_out_to_Subtract13_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Subtract13_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Subtract13_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Subtract13_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Subtract13_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No216_out_to_Add56_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No217_out_to_Add56_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Add56_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Add56_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Add56_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Add56_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No218_out_to_Product43_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No219_out_to_Product43_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Product43_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Product43_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product43_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product43_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No220_out_to_Product115_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No221_out_to_Product115_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Product115_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Product115_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product115_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out_to_MUX_Product115_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No222_out_to_Product214_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No223_out_to_Product214_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Product214_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Product214_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product214_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product214_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No224_out_to_Product314_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No225_out_to_Product314_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product314_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out_to_MUX_Product314_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Product314_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Product314_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No226_out_to_Subtract15_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No227_out_to_Subtract15_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Subtract15_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Subtract15_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Subtract15_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Subtract15_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No228_out_to_Add57_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No229_out_to_Add57_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Add57_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Add57_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Add57_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Add57_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No230_out_to_Product44_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No231_out_to_Product44_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Product44_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Product44_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Product44_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Product44_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No232_out_to_Product116_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No233_out_to_Product116_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Product116_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Product116_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Product116_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Product116_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No234_out_to_Product215_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No235_out_to_Product215_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Product215_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Product215_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Product215_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Product215_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No236_out_to_Product315_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No237_out_to_Product315_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Product315_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Product315_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Product315_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Product315_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No238_out_to_Subtract16_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No239_out_to_Subtract16_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Subtract16_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Subtract16_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Subtract16_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Subtract16_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No240_out_to_Add58_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No241_out_to_Add58_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Add58_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Add58_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Add58_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Add58_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No242_out_to_Product45_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No243_out_to_Product45_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Product45_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Product45_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out_to_MUX_Product45_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Product45_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No244_out_to_Product117_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No245_out_to_Product117_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Product117_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Product117_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Product117_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Product117_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No246_out_to_Product216_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No247_out_to_Product216_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Product216_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Product216_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out_to_MUX_Product216_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Product216_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No248_out_to_Product316_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No249_out_to_Product316_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Product316_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Product316_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Product316_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Product316_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No250_out_to_Subtract17_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No251_out_to_Subtract17_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No252_out_to_Add59_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No253_out_to_Add59_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Add59_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Add59_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Add59_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Add59_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No254_out_to_Product46_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No255_out_to_Product46_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Product46_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Product46_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out_to_MUX_Product46_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Product46_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No256_out_to_Product118_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No257_out_to_Product118_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Product118_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Product118_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Product118_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Product118_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No258_out_to_Product217_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No259_out_to_Product217_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Product217_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Product217_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out_to_MUX_Product217_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Product217_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No260_out_to_Product317_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No261_out_to_Product317_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Product317_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Product317_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Product317_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Product317_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No262_out_to_Subtract18_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No263_out_to_Subtract18_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Subtract18_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Subtract18_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Subtract18_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Subtract18_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No264_out_to_Add61_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No265_out_to_Add61_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Add61_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Add61_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Add61_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Add61_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No266_out_to_Product48_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No267_out_to_Product48_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Product48_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out_to_MUX_Product48_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product48_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product48_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No268_out_to_Product120_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No269_out_to_Product120_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Product120_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out_to_MUX_Product120_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product120_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Product120_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No270_out_to_Product219_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No271_out_to_Product219_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Product219_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Product219_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product219_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product219_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No272_out_to_Product319_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No273_out_to_Product319_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product319_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Product319_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Product319_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Product319_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No274_out_to_Subtract20_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No275_out_to_Subtract20_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No276_out_to_Add63_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No277_out_to_Add63_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Add63_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Add63_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Add63_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Add63_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No278_out_to_Product50_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No279_out_to_Product50_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Product50_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out_to_MUX_Product50_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Product50_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Product50_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No280_out_to_Product122_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No281_out_to_Product122_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Product122_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out_to_MUX_Product122_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Product122_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product122_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No282_out_to_Product221_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No283_out_to_Product221_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Product221_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out_to_MUX_Product221_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Product221_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Product221_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No284_out_to_Product321_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No285_out_to_Product321_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Product321_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product321_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Product321_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out_to_MUX_Product321_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No286_out_to_Subtract22_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No287_out_to_Subtract22_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Subtract22_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Subtract22_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Subtract22_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Subtract22_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No288_out_to_Add65_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No289_out_to_Add65_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Add65_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out_to_MUX_Add65_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Add65_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Add65_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No290_out_to_Product52_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No291_out_to_Product52_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Product52_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Product52_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Product52_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Product52_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No292_out_to_Product124_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No293_out_to_Product124_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Product124_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Product124_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Product124_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out_to_MUX_Product124_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No294_out_to_Product223_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No295_out_to_Product223_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Product223_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Product223_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Product223_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Product223_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No296_out_to_Product323_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No297_out_to_Product323_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Product323_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out_to_MUX_Product323_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Product323_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Product323_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No298_out_to_Subtract24_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No299_out_to_Subtract24_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Subtract24_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Subtract24_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Subtract24_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Subtract24_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No300_out_to_Add66_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No301_out_to_Add66_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out_to_MUX_Add66_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Add66_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Add66_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Add66_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No302_out_to_Product53_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No303_out_to_Product53_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Product53_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Product53_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product53_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product53_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No304_out_to_Product125_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No305_out_to_Product125_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Product125_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Product125_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product125_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Product125_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No306_out_to_Product224_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No307_out_to_Product224_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Product224_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Product224_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product224_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product224_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No308_out_to_Product324_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No309_out_to_Product324_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product324_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Product324_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Product324_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Product324_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No310_out_to_Subtract25_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No311_out_to_Subtract25_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Subtract25_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Subtract25_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Subtract25_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Subtract25_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No312_out_to_Add67_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No313_out_to_Add67_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Add67_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Add67_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Add67_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Add67_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No314_out_to_Product54_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No315_out_to_Product54_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Product54_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Product54_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Product54_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Product54_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No316_out_to_Product126_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No317_out_to_Product126_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Product126_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Product126_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Product126_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Product126_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No318_out_to_Product225_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No319_out_to_Product225_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Product225_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Product225_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Product225_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Product225_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No320_out_to_Product325_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No321_out_to_Product325_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Product325_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Product325_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Product325_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Product325_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No322_out_to_Subtract26_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No323_out_to_Subtract26_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Subtract26_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Subtract26_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Subtract26_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Subtract26_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No324_out_to_Add68_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No325_out_to_Add68_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Add68_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Add68_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Add68_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Add68_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No326_out_to_Product55_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No327_out_to_Product55_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Product55_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out_to_MUX_Product55_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Product55_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Product55_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No328_out_to_Product127_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No329_out_to_Product127_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Product127_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out_to_MUX_Product127_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Product127_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Product127_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No330_out_to_Product226_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No331_out_to_Product226_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Product226_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out_to_MUX_Product226_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Product226_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Product226_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No332_out_to_Product326_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No333_out_to_Product326_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Product326_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Product326_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Product326_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out_to_MUX_Product326_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No334_out_to_Subtract27_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No335_out_to_Subtract27_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Subtract27_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Subtract27_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Subtract27_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Subtract27_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No336_out_to_Add83_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No337_out_to_Add83_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Add83_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Add83_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Add83_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Add83_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No338_out_to_Product70_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No339_out_to_Product70_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Product70_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Product70_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product70_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product70_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No340_out_to_Product142_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No341_out_to_Product142_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Product142_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Product142_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Product142_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product142_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No342_out_to_Product241_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No343_out_to_Product241_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Product241_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Product241_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product241_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product241_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No344_out_to_Product341_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No345_out_to_Product341_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Product341_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product341_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Product341_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Product341_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No346_out_to_Subtract42_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No347_out_to_Subtract42_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Subtract42_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Subtract42_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Subtract42_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Subtract42_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No348_out_to_Add84_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No349_out_to_Add84_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out_to_MUX_Add84_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out_to_MUX_Add84_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Add84_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Add84_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No350_out_to_Product71_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No351_out_to_Product71_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Product71_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Product71_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product71_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Product71_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No352_out_to_Product143_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No353_out_to_Product143_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Product143_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Product143_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product143_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Product143_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No354_out_to_Product242_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No355_out_to_Product242_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Product242_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Product242_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product242_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Product242_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No356_out_to_Product342_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No357_out_to_Product342_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product342_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Product342_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Product342_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Product342_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No358_out_to_Subtract43_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No359_out_to_Subtract43_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Subtract43_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Subtract43_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Subtract43_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Subtract43_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No360_out_to_Add85_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No361_out_to_Add85_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Add85_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Add85_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Add85_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Add85_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No362_out_to_Product72_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No363_out_to_Product72_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Product72_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Product72_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Product72_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Product72_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No364_out_to_Product144_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No365_out_to_Product144_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Product144_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Product144_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Product144_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Product144_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No366_out_to_Product243_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No367_out_to_Product243_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Product243_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Product243_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Product243_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Product243_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No368_out_to_Product343_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No369_out_to_Product343_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Product343_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Product343_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Product343_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Product343_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No370_out_to_Subtract44_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No371_out_to_Subtract44_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Subtract44_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Subtract44_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Subtract44_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Subtract44_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No372_out_to_Subtract45_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No373_out_to_Subtract45_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Subtract45_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract45_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Subtract45_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract45_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No374_out_to_Add87_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No375_out_to_Add87_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out_to_MUX_Add87_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out_to_MUX_Add87_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Add87_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Add87_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No376_out_to_Product74_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No377_out_to_Product74_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Product74_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Product74_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Product74_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product74_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No378_out_to_Product146_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No379_out_to_Product146_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Product146_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Product146_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Product146_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product146_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No380_out_to_Product245_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No381_out_to_Product245_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Product245_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Product245_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Product245_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product245_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No382_out_to_Product345_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No383_out_to_Product345_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Product345_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product345_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Product345_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Product345_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No384_out_to_Subtract46_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No385_out_to_Subtract46_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Subtract46_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Subtract46_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Subtract46_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out_to_MUX_Subtract46_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No386_out_to_Subtract47_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No387_out_to_Subtract47_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Subtract47_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract47_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Subtract47_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract47_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No388_out_to_Subtract48_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No389_out_to_Subtract48_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Subtract48_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract48_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Subtract48_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract48_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No390_out_to_Subtract49_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No391_out_to_Subtract49_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Subtract49_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Subtract49_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out_to_MUX_Subtract49_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Subtract49_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No392_out_to_Subtract50_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No393_out_to_Subtract50_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Subtract50_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract50_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Subtract50_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract50_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No394_out_to_Subtract52_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No395_out_to_Subtract52_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Subtract52_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Subtract52_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Subtract52_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Subtract52_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No396_out_to_Subtract112_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No397_out_to_Subtract112_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Subtract112_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Subtract112_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Subtract112_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Subtract112_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No398_out_to_Subtract114_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No399_out_to_Subtract114_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Subtract114_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Subtract114_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Subtract114_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Subtract114_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No400_out_to_Subtract55_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No401_out_to_Subtract55_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Subtract55_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Subtract55_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Subtract55_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Subtract55_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No402_out_to_Subtract115_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No403_out_to_Subtract115_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Subtract115_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Subtract115_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Subtract115_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Subtract115_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No404_out_to_Subtract56_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No405_out_to_Subtract56_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Subtract56_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Subtract56_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Subtract56_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Subtract56_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No406_out_to_Subtract116_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No407_out_to_Subtract116_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No49_out_to_MUX_Subtract116_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Subtract116_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No51_out_to_MUX_Subtract116_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Subtract116_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No408_out_to_Subtract57_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No409_out_to_Subtract57_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No48_out_to_MUX_Subtract57_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Subtract57_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No50_out_to_MUX_Subtract57_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Subtract57_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No410_out_to_Subtract117_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No411_out_to_Subtract117_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No41_out_to_MUX_Subtract117_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Subtract117_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No43_out_to_MUX_Subtract117_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Subtract117_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No412_out_to_Subtract59_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No413_out_to_Subtract59_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No40_out_to_MUX_Subtract59_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Subtract59_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No42_out_to_MUX_Subtract59_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Subtract59_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No414_out_to_Subtract119_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No415_out_to_Subtract119_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No45_out_to_MUX_Subtract119_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Subtract119_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No53_out_to_MUX_Subtract119_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Subtract119_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No416_out_to_Subtract62_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No417_out_to_Subtract62_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No44_out_to_MUX_Subtract62_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract62_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No52_out_to_MUX_Subtract62_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract62_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No418_out_to_Subtract122_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No419_out_to_Subtract122_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No47_out_to_MUX_Subtract122_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Subtract122_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No55_out_to_MUX_Subtract122_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract122_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No420_out_to_Subtract63_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No421_out_to_Subtract63_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No46_out_to_MUX_Subtract63_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Subtract63_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No54_out_to_MUX_Subtract63_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Subtract63_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No422_out_to_Subtract123_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No423_out_to_Subtract123_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Subtract123_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Subtract123_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Subtract123_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Subtract123_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No424_out_to_Subtract127_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No425_out_to_Subtract127_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Subtract127_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract127_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Subtract127_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract127_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No426_out_to_Subtract68_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No427_out_to_Subtract68_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Subtract68_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract68_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Subtract68_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Subtract68_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No428_out_to_Subtract71_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No429_out_to_Subtract71_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Subtract71_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract71_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Subtract71_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract71_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No430_out_to_Subtract131_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No431_out_to_Subtract131_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Subtract131_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract131_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Subtract131_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract131_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No432_out_to_Subtract72_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No433_out_to_Subtract72_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Subtract72_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract72_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Subtract72_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract72_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No434_out_to_Subtract132_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No435_out_to_Subtract132_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Subtract132_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract132_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Subtract132_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract132_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No436_out_to_Subtract74_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No437_out_to_Subtract74_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Subtract74_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract74_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out_to_MUX_Subtract74_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract74_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No438_out_to_Subtract134_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No439_out_to_Subtract134_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Subtract134_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract134_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out_to_MUX_Subtract134_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract134_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No440_out_to_Subtract75_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No441_out_to_Subtract75_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out_to_MUX_Subtract75_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract75_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Subtract75_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract75_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No442_out_to_Subtract135_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No443_out_to_Subtract135_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Subtract135_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Subtract135_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Subtract135_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract135_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No444_out_to_Subtract80_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No445_out_to_Subtract80_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Subtract80_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Subtract80_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Subtract80_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Subtract80_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No446_out_to_Subtract140_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No447_out_to_Subtract140_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Subtract140_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Subtract140_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Subtract140_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out_to_MUX_Subtract140_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   ModCount21_instance: ModuloCounter_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Counter_out => ModCount21_out);
x0_re_IEEE <= x0_re;
   x0_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x0_re_out,
                 X => x0_re_IEEE);
x0_im_IEEE <= x0_im;
   x0_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x0_im_out,
                 X => x0_im_IEEE);
x1_re_IEEE <= x1_re;
   x1_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x1_re_out,
                 X => x1_re_IEEE);
x1_im_IEEE <= x1_im;
   x1_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x1_im_out,
                 X => x1_im_IEEE);
x2_re_IEEE <= x2_re;
   x2_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x2_re_out,
                 X => x2_re_IEEE);
x2_im_IEEE <= x2_im;
   x2_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x2_im_out,
                 X => x2_im_IEEE);
x3_re_IEEE <= x3_re;
   x3_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x3_re_out,
                 X => x3_re_IEEE);
x3_im_IEEE <= x3_im;
   x3_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x3_im_out,
                 X => x3_im_IEEE);
x4_re_IEEE <= x4_re;
   x4_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x4_re_out,
                 X => x4_re_IEEE);
x4_im_IEEE <= x4_im;
   x4_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x4_im_out,
                 X => x4_im_IEEE);
x5_re_IEEE <= x5_re;
   x5_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x5_re_out,
                 X => x5_re_IEEE);
x5_im_IEEE <= x5_im;
   x5_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x5_im_out,
                 X => x5_im_IEEE);
x6_re_IEEE <= x6_re;
   x6_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x6_re_out,
                 X => x6_re_IEEE);
x6_im_IEEE <= x6_im;
   x6_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x6_im_out,
                 X => x6_im_IEEE);
x7_re_IEEE <= x7_re;
   x7_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x7_re_out,
                 X => x7_re_IEEE);
x7_im_IEEE <= x7_im;
   x7_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x7_im_out,
                 X => x7_im_IEEE);
x8_re_IEEE <= x8_re;
   x8_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x8_re_out,
                 X => x8_re_IEEE);
x8_im_IEEE <= x8_im;
   x8_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x8_im_out,
                 X => x8_im_IEEE);
x9_re_IEEE <= x9_re;
   x9_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x9_re_out,
                 X => x9_re_IEEE);
x9_im_IEEE <= x9_im;
   x9_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x9_im_out,
                 X => x9_im_IEEE);
x10_re_IEEE <= x10_re;
   x10_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x10_re_out,
                 X => x10_re_IEEE);
x10_im_IEEE <= x10_im;
   x10_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x10_im_out,
                 X => x10_im_IEEE);
x11_re_IEEE <= x11_re;
   x11_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x11_re_out,
                 X => x11_re_IEEE);
x11_im_IEEE <= x11_im;
   x11_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x11_im_out,
                 X => x11_im_IEEE);
x12_re_IEEE <= x12_re;
   x12_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x12_re_out,
                 X => x12_re_IEEE);
x12_im_IEEE <= x12_im;
   x12_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x12_im_out,
                 X => x12_im_IEEE);
x13_re_IEEE <= x13_re;
   x13_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x13_re_out,
                 X => x13_re_IEEE);
x13_im_IEEE <= x13_im;
   x13_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x13_im_out,
                 X => x13_im_IEEE);
x14_re_IEEE <= x14_re;
   x14_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x14_re_out,
                 X => x14_re_IEEE);
x14_im_IEEE <= x14_im;
   x14_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x14_im_out,
                 X => x14_im_IEEE);
x15_re_IEEE <= x15_re;
   x15_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x15_re_out,
                 X => x15_re_IEEE);
x15_im_IEEE <= x15_im;
   x15_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x15_im_out,
                 X => x15_im_IEEE);
   y0_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y0_re_IEEE,
                 X => Delay1No_out);
y0_re <= y0_re_IEEE;

   Delay1No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg42_out,
                 Y => Delay1No_out);
   y0_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y0_im_IEEE,
                 X => Delay1No1_out);
y0_im <= y0_im_IEEE;

   Delay1No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg43_out,
                 Y => Delay1No1_out);
   y1_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y1_re_IEEE,
                 X => Delay1No2_out);
y1_re <= y1_re_IEEE;

   Delay1No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg56_out,
                 Y => Delay1No2_out);
   y1_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y1_im_IEEE,
                 X => Delay1No3_out);
y1_im <= y1_im_IEEE;

   Delay1No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg58_out,
                 Y => Delay1No3_out);
   y2_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y2_re_IEEE,
                 X => Delay1No4_out);
y2_re <= y2_re_IEEE;

   Delay1No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg48_out,
                 Y => Delay1No4_out);
   y2_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y2_im_IEEE,
                 X => Delay1No5_out);
y2_im <= y2_im_IEEE;

   Delay1No5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg50_out,
                 Y => Delay1No5_out);
   y3_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y3_re_IEEE,
                 X => Delay1No6_out);
y3_re <= y3_re_IEEE;

   Delay1No6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg66_out,
                 Y => Delay1No6_out);
   y3_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y3_im_IEEE,
                 X => Delay1No7_out);
y3_im <= y3_im_IEEE;

   Delay1No7_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg68_out,
                 Y => Delay1No7_out);
   y4_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y4_re_IEEE,
                 X => Delay1No8_out);
y4_re <= y4_re_IEEE;

   Delay1No8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg44_out,
                 Y => Delay1No8_out);
   y4_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y4_im_IEEE,
                 X => Delay1No9_out);
y4_im <= y4_im_IEEE;

   Delay1No9_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg46_out,
                 Y => Delay1No9_out);
   y5_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y5_re_IEEE,
                 X => Delay1No10_out);
y5_re <= y5_re_IEEE;

   Delay1No10_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg60_out,
                 Y => Delay1No10_out);
   y5_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y5_im_IEEE,
                 X => Delay1No11_out);
y5_im <= y5_im_IEEE;

   Delay1No11_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg62_out,
                 Y => Delay1No11_out);
   y6_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y6_re_IEEE,
                 X => Delay1No12_out);
y6_re <= y6_re_IEEE;

   Delay1No12_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg52_out,
                 Y => Delay1No12_out);
   y6_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y6_im_IEEE,
                 X => Delay1No13_out);
y6_im <= y6_im_IEEE;

   Delay1No13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg54_out,
                 Y => Delay1No13_out);
   y7_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y7_re_IEEE,
                 X => Delay1No14_out);
y7_re <= y7_re_IEEE;

   Delay1No14_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg69_out,
                 Y => Delay1No14_out);
   y7_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y7_im_IEEE,
                 X => Delay1No15_out);
y7_im <= y7_im_IEEE;

   Delay1No15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg70_out,
                 Y => Delay1No15_out);
   y8_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y8_re_IEEE,
                 X => Delay1No16_out);
y8_re <= y8_re_IEEE;

   Delay1No16_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg242_out,
                 Y => Delay1No16_out);
   y8_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y8_im_IEEE,
                 X => Delay1No17_out);
y8_im <= y8_im_IEEE;

   Delay1No17_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg244_out,
                 Y => Delay1No17_out);
   y9_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y9_re_IEEE,
                 X => Delay1No18_out);
y9_re <= y9_re_IEEE;

   Delay1No18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg246_out,
                 Y => Delay1No18_out);
   y9_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y9_im_IEEE,
                 X => Delay1No19_out);
y9_im <= y9_im_IEEE;

   Delay1No19_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg247_out,
                 Y => Delay1No19_out);
   y10_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y10_re_IEEE,
                 X => Delay1No20_out);
y10_re <= y10_re_IEEE;

   Delay1No20_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg207_out,
                 Y => Delay1No20_out);
   y10_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y10_im_IEEE,
                 X => Delay1No21_out);
y10_im <= y10_im_IEEE;

   Delay1No21_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg213_out,
                 Y => Delay1No21_out);
   y11_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y11_re_IEEE,
                 X => Delay1No22_out);
y11_re <= y11_re_IEEE;

   Delay1No22_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg250_out,
                 Y => Delay1No22_out);
   y11_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y11_im_IEEE,
                 X => Delay1No23_out);
y11_im <= y11_im_IEEE;

   Delay1No23_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg251_out,
                 Y => Delay1No23_out);
   y12_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y12_re_IEEE,
                 X => Delay1No24_out);
y12_re <= y12_re_IEEE;

   Delay1No24_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg245_out,
                 Y => Delay1No24_out);
   y12_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y12_im_IEEE,
                 X => Delay1No25_out);
y12_im <= y12_im_IEEE;

   Delay1No25_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg201_out,
                 Y => Delay1No25_out);
   y13_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y13_re_IEEE,
                 X => Delay1No26_out);
y13_re <= y13_re_IEEE;

   Delay1No26_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg248_out,
                 Y => Delay1No26_out);
   y13_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y13_im_IEEE,
                 X => Delay1No27_out);
y13_im <= y13_im_IEEE;

   Delay1No27_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg249_out,
                 Y => Delay1No27_out);
   y14_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y14_re_IEEE,
                 X => Delay1No28_out);
y14_re <= y14_re_IEEE;

   Delay1No28_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg220_out,
                 Y => Delay1No28_out);
   y14_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y14_im_IEEE,
                 X => Delay1No29_out);
y14_im <= y14_im_IEEE;

   Delay1No29_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg224_out,
                 Y => Delay1No29_out);
   y15_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y15_re_IEEE,
                 X => Delay1No30_out);
y15_re <= y15_re_IEEE;

   Delay1No30_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg252_out,
                 Y => Delay1No30_out);
   y15_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y15_im_IEEE,
                 X => Delay1No31_out);
y15_im <= y15_im_IEEE;

   Delay1No31_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg253_out,
                 Y => Delay1No31_out);

Delay1No32_out_to_Add2_impl_parent_implementedSystem_port_0_cast <= Delay1No32_out;
Delay1No33_out_to_Add2_impl_parent_implementedSystem_port_1_cast <= Delay1No33_out;
   Add2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_impl_out,
                 X => Delay1No32_out_to_Add2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No33_out_to_Add2_impl_parent_implementedSystem_port_1_cast);

Delay2No_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_1_cast <= Delay2No_out;
SharedReg84_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg84_out;
   MUX_Add2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg84_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add2_impl_0_out);

   Delay1No32_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_impl_0_out,
                 Y => Delay1No32_out);

Delay2No8_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_1_cast <= Delay2No8_out;
SharedReg106_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg106_out;
   MUX_Add2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No8_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg106_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add2_impl_1_out);

   Delay1No33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_impl_1_out,
                 Y => Delay1No33_out);

Delay1No34_out_to_Add11_impl_parent_implementedSystem_port_0_cast <= Delay1No34_out;
Delay1No35_out_to_Add11_impl_parent_implementedSystem_port_1_cast <= Delay1No35_out;
   Add11_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_impl_out,
                 X => Delay1No34_out_to_Add11_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No35_out_to_Add11_impl_parent_implementedSystem_port_1_cast);

Delay2No1_out_to_MUX_Add11_impl_0_parent_implementedSystem_port_1_cast <= Delay2No1_out;
SharedReg2_out_to_MUX_Add11_impl_0_parent_implementedSystem_port_2_cast <= SharedReg2_out;
   MUX_Add11_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No1_out_to_MUX_Add11_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg2_out_to_MUX_Add11_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add11_impl_0_out);

   Delay1No34_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_impl_0_out,
                 Y => Delay1No34_out);

Delay2No9_out_to_MUX_Add11_impl_1_parent_implementedSystem_port_1_cast <= Delay2No9_out;
SharedReg18_out_to_MUX_Add11_impl_1_parent_implementedSystem_port_2_cast <= SharedReg18_out;
   MUX_Add11_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No9_out_to_MUX_Add11_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg18_out_to_MUX_Add11_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add11_impl_1_out);

   Delay1No35_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_impl_1_out,
                 Y => Delay1No35_out);

Delay1No36_out_to_Add12_impl_parent_implementedSystem_port_0_cast <= Delay1No36_out;
Delay1No37_out_to_Add12_impl_parent_implementedSystem_port_1_cast <= Delay1No37_out;
   Add12_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add12_impl_out,
                 X => Delay1No36_out_to_Add12_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No37_out_to_Add12_impl_parent_implementedSystem_port_1_cast);

SharedReg89_out_to_MUX_Add12_impl_0_parent_implementedSystem_port_1_cast <= SharedReg89_out;
SharedReg3_out_to_MUX_Add12_impl_0_parent_implementedSystem_port_2_cast <= SharedReg3_out;
   MUX_Add12_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg89_out_to_MUX_Add12_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg3_out_to_MUX_Add12_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add12_impl_0_out);

   Delay1No36_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_impl_0_out,
                 Y => Delay1No36_out);

SharedReg220_out_to_MUX_Add12_impl_1_parent_implementedSystem_port_1_cast <= SharedReg220_out;
SharedReg19_out_to_MUX_Add12_impl_1_parent_implementedSystem_port_2_cast <= SharedReg19_out;
   MUX_Add12_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg220_out_to_MUX_Add12_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg19_out_to_MUX_Add12_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add12_impl_1_out);

   Delay1No37_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_impl_1_out,
                 Y => Delay1No37_out);

Delay1No38_out_to_Add13_impl_parent_implementedSystem_port_0_cast <= Delay1No38_out;
Delay1No39_out_to_Add13_impl_parent_implementedSystem_port_1_cast <= Delay1No39_out;
   Add13_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add13_impl_out,
                 X => Delay1No38_out_to_Add13_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No39_out_to_Add13_impl_parent_implementedSystem_port_1_cast);

SharedReg90_out_to_MUX_Add13_impl_0_parent_implementedSystem_port_1_cast <= SharedReg90_out;
SharedReg183_out_to_MUX_Add13_impl_0_parent_implementedSystem_port_2_cast <= SharedReg183_out;
   MUX_Add13_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg90_out_to_MUX_Add13_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg183_out_to_MUX_Add13_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add13_impl_0_out);

   Delay1No38_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add13_impl_0_out,
                 Y => Delay1No38_out);

SharedReg215_out_to_MUX_Add13_impl_1_parent_implementedSystem_port_1_cast <= SharedReg215_out;
SharedReg221_out_to_MUX_Add13_impl_1_parent_implementedSystem_port_2_cast <= SharedReg221_out;
   MUX_Add13_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg215_out_to_MUX_Add13_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg221_out_to_MUX_Add13_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add13_impl_1_out);

   Delay1No39_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add13_impl_1_out,
                 Y => Delay1No39_out);

Delay1No40_out_to_Add14_impl_parent_implementedSystem_port_0_cast <= Delay1No40_out;
Delay1No41_out_to_Add14_impl_parent_implementedSystem_port_1_cast <= Delay1No41_out;
   Add14_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add14_impl_out,
                 X => Delay1No40_out_to_Add14_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No41_out_to_Add14_impl_parent_implementedSystem_port_1_cast);

SharedReg83_out_to_MUX_Add14_impl_0_parent_implementedSystem_port_1_cast <= SharedReg83_out;
SharedReg178_out_to_MUX_Add14_impl_0_parent_implementedSystem_port_2_cast <= SharedReg178_out;
   MUX_Add14_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg83_out_to_MUX_Add14_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg178_out_to_MUX_Add14_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add14_impl_0_out);

   Delay1No40_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add14_impl_0_out,
                 Y => Delay1No40_out);

SharedReg123_out_to_MUX_Add14_impl_1_parent_implementedSystem_port_1_cast <= SharedReg123_out;
SharedReg202_out_to_MUX_Add14_impl_1_parent_implementedSystem_port_2_cast <= SharedReg202_out;
   MUX_Add14_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg123_out_to_MUX_Add14_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg202_out_to_MUX_Add14_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add14_impl_1_out);

   Delay1No41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add14_impl_1_out,
                 Y => Delay1No41_out);

Delay1No42_out_to_Add6_impl_parent_implementedSystem_port_0_cast <= Delay1No42_out;
Delay1No43_out_to_Add6_impl_parent_implementedSystem_port_1_cast <= Delay1No43_out;
   Add6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add6_impl_out,
                 X => Delay1No42_out_to_Add6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No43_out_to_Add6_impl_parent_implementedSystem_port_1_cast);

SharedReg84_out_to_MUX_Add6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg84_out;
SharedReg222_out_to_MUX_Add6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg222_out;
   MUX_Add6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg84_out_to_MUX_Add6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg222_out_to_MUX_Add6_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add6_impl_0_out);

   Delay1No42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add6_impl_0_out,
                 Y => Delay1No42_out);

SharedReg124_out_to_MUX_Add6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg124_out;
SharedReg99_out_to_MUX_Add6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg99_out;
   MUX_Add6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg124_out_to_MUX_Add6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg99_out_to_MUX_Add6_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add6_impl_1_out);

   Delay1No43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add6_impl_1_out,
                 Y => Delay1No43_out);

Delay1No44_out_to_Add15_impl_parent_implementedSystem_port_0_cast <= Delay1No44_out;
Delay1No45_out_to_Add15_impl_parent_implementedSystem_port_1_cast <= Delay1No45_out;
   Add15_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add15_impl_out,
                 X => Delay1No44_out_to_Add15_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No45_out_to_Add15_impl_parent_implementedSystem_port_1_cast);

SharedReg99_out_to_MUX_Add15_impl_0_parent_implementedSystem_port_1_cast <= SharedReg99_out;
SharedReg208_out_to_MUX_Add15_impl_0_parent_implementedSystem_port_2_cast <= SharedReg208_out;
   MUX_Add15_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg99_out_to_MUX_Add15_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg208_out_to_MUX_Add15_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add15_impl_0_out);

   Delay1No44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add15_impl_0_out,
                 Y => Delay1No44_out);

SharedReg105_out_to_MUX_Add15_impl_1_parent_implementedSystem_port_1_cast <= SharedReg105_out;
SharedReg94_out_to_MUX_Add15_impl_1_parent_implementedSystem_port_2_cast <= SharedReg94_out;
   MUX_Add15_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg105_out_to_MUX_Add15_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg94_out_to_MUX_Add15_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add15_impl_1_out);

   Delay1No45_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add15_impl_1_out,
                 Y => Delay1No45_out);

Delay1No46_out_to_Add7_impl_parent_implementedSystem_port_0_cast <= Delay1No46_out;
Delay1No47_out_to_Add7_impl_parent_implementedSystem_port_1_cast <= Delay1No47_out;
   Add7_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add7_impl_out,
                 X => Delay1No46_out_to_Add7_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No47_out_to_Add7_impl_parent_implementedSystem_port_1_cast);

SharedReg94_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_1_cast <= SharedReg94_out;
SharedReg223_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_2_cast <= SharedReg223_out;
   MUX_Add7_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg94_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg223_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add7_impl_0_out);

   Delay1No46_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add7_impl_0_out,
                 Y => Delay1No46_out);

SharedReg100_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_1_cast <= SharedReg100_out;
SharedReg105_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_2_cast <= SharedReg105_out;
   MUX_Add7_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg100_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg105_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add7_impl_1_out);

   Delay1No47_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add7_impl_1_out,
                 Y => Delay1No47_out);

Delay1No48_out_to_Add16_impl_parent_implementedSystem_port_0_cast <= Delay1No48_out;
Delay1No49_out_to_Add16_impl_parent_implementedSystem_port_1_cast <= Delay1No49_out;
   Add16_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add16_impl_out,
                 X => Delay1No48_out_to_Add16_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No49_out_to_Add16_impl_parent_implementedSystem_port_1_cast);

Delay2No2_out_to_MUX_Add16_impl_0_parent_implementedSystem_port_1_cast <= Delay2No2_out;
SharedReg215_out_to_MUX_Add16_impl_0_parent_implementedSystem_port_2_cast <= SharedReg215_out;
   MUX_Add16_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No2_out_to_MUX_Add16_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg215_out_to_MUX_Add16_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add16_impl_0_out);

   Delay1No48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add16_impl_0_out,
                 Y => Delay1No48_out);

Delay2No10_out_to_MUX_Add16_impl_1_parent_implementedSystem_port_1_cast <= Delay2No10_out;
SharedReg100_out_to_MUX_Add16_impl_1_parent_implementedSystem_port_2_cast <= SharedReg100_out;
   MUX_Add16_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No10_out_to_MUX_Add16_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg100_out_to_MUX_Add16_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add16_impl_1_out);

   Delay1No49_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add16_impl_1_out,
                 Y => Delay1No49_out);

Delay1No50_out_to_Add8_impl_parent_implementedSystem_port_0_cast <= Delay1No50_out;
Delay1No51_out_to_Add8_impl_parent_implementedSystem_port_1_cast <= Delay1No51_out;
   Add8_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add8_impl_out,
                 X => Delay1No50_out_to_Add8_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No51_out_to_Add8_impl_parent_implementedSystem_port_1_cast);

Delay2No3_out_to_MUX_Add8_impl_0_parent_implementedSystem_port_1_cast <= Delay2No3_out;
SharedReg89_out_to_MUX_Add8_impl_0_parent_implementedSystem_port_2_cast <= SharedReg89_out;
   MUX_Add8_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No3_out_to_MUX_Add8_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg89_out_to_MUX_Add8_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add8_impl_0_out);

   Delay1No50_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add8_impl_0_out,
                 Y => Delay1No50_out);

Delay2No11_out_to_MUX_Add8_impl_1_parent_implementedSystem_port_1_cast <= Delay2No11_out;
SharedReg111_out_to_MUX_Add8_impl_1_parent_implementedSystem_port_2_cast <= SharedReg111_out;
   MUX_Add8_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No11_out_to_MUX_Add8_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg111_out_to_MUX_Add8_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add8_impl_1_out);

   Delay1No51_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add8_impl_1_out,
                 Y => Delay1No51_out);

Delay1No52_out_to_Add9_impl_parent_implementedSystem_port_0_cast <= Delay1No52_out;
Delay1No53_out_to_Add9_impl_parent_implementedSystem_port_1_cast <= Delay1No53_out;
   Add9_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add9_impl_out,
                 X => Delay1No52_out_to_Add9_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No53_out_to_Add9_impl_parent_implementedSystem_port_1_cast);

SharedReg111_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_1_cast <= SharedReg111_out;
SharedReg81_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_2_cast <= SharedReg81_out;
   MUX_Add9_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg111_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg81_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add9_impl_0_out);

   Delay1No52_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add9_impl_0_out,
                 Y => Delay1No52_out);

SharedReg117_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_1_cast <= SharedReg117_out;
SharedReg117_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_2_cast <= SharedReg117_out;
   MUX_Add9_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg117_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg117_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add9_impl_1_out);

   Delay1No53_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add9_impl_1_out,
                 Y => Delay1No53_out);

Delay1No54_out_to_Add18_impl_parent_implementedSystem_port_0_cast <= Delay1No54_out;
Delay1No55_out_to_Add18_impl_parent_implementedSystem_port_1_cast <= Delay1No55_out;
   Add18_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add18_impl_out,
                 X => Delay1No54_out_to_Add18_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No55_out_to_Add18_impl_parent_implementedSystem_port_1_cast);

SharedReg106_out_to_MUX_Add18_impl_0_parent_implementedSystem_port_1_cast <= SharedReg106_out;
SharedReg90_out_to_MUX_Add18_impl_0_parent_implementedSystem_port_2_cast <= SharedReg90_out;
   MUX_Add18_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg106_out_to_MUX_Add18_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg90_out_to_MUX_Add18_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add18_impl_0_out);

   Delay1No54_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add18_impl_0_out,
                 Y => Delay1No54_out);

SharedReg112_out_to_MUX_Add18_impl_1_parent_implementedSystem_port_1_cast <= SharedReg112_out;
SharedReg112_out_to_MUX_Add18_impl_1_parent_implementedSystem_port_2_cast <= SharedReg112_out;
   MUX_Add18_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg112_out_to_MUX_Add18_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg112_out_to_MUX_Add18_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add18_impl_1_out);

   Delay1No55_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add18_impl_1_out,
                 Y => Delay1No55_out);

Delay1No56_out_to_Add20_impl_parent_implementedSystem_port_0_cast <= Delay1No56_out;
Delay1No57_out_to_Add20_impl_parent_implementedSystem_port_1_cast <= Delay1No57_out;
   Add20_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add20_impl_out,
                 X => Delay1No56_out_to_Add20_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No57_out_to_Add20_impl_parent_implementedSystem_port_1_cast);

SharedReg171_out_to_MUX_Add20_impl_0_parent_implementedSystem_port_1_cast <= SharedReg171_out;
SharedReg123_out_to_MUX_Add20_impl_0_parent_implementedSystem_port_2_cast <= SharedReg123_out;
   MUX_Add20_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg171_out_to_MUX_Add20_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg123_out_to_MUX_Add20_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add20_impl_0_out);

   Delay1No56_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add20_impl_0_out,
                 Y => Delay1No56_out);

SharedReg177_out_to_MUX_Add20_impl_1_parent_implementedSystem_port_1_cast <= SharedReg177_out;
SharedReg165_out_to_MUX_Add20_impl_1_parent_implementedSystem_port_2_cast <= SharedReg165_out;
   MUX_Add20_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg177_out_to_MUX_Add20_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg165_out_to_MUX_Add20_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add20_impl_1_out);

   Delay1No57_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add20_impl_1_out,
                 Y => Delay1No57_out);

Delay1No58_out_to_Add110_impl_parent_implementedSystem_port_0_cast <= Delay1No58_out;
Delay1No59_out_to_Add110_impl_parent_implementedSystem_port_1_cast <= Delay1No59_out;
   Add110_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add110_impl_out,
                 X => Delay1No58_out_to_Add110_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No59_out_to_Add110_impl_parent_implementedSystem_port_1_cast);

SharedReg166_out_to_MUX_Add110_impl_0_parent_implementedSystem_port_1_cast <= SharedReg166_out;
SharedReg118_out_to_MUX_Add110_impl_0_parent_implementedSystem_port_2_cast <= SharedReg118_out;
   MUX_Add110_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg166_out_to_MUX_Add110_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg118_out_to_MUX_Add110_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add110_impl_0_out);

   Delay1No58_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add110_impl_0_out,
                 Y => Delay1No58_out);

SharedReg172_out_to_MUX_Add110_impl_1_parent_implementedSystem_port_1_cast <= SharedReg172_out;
SharedReg160_out_to_MUX_Add110_impl_1_parent_implementedSystem_port_2_cast <= SharedReg160_out;
   MUX_Add110_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg172_out_to_MUX_Add110_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg160_out_to_MUX_Add110_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add110_impl_1_out);

   Delay1No59_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add110_impl_1_out,
                 Y => Delay1No59_out);

Delay1No60_out_to_Add22_impl_parent_implementedSystem_port_0_cast <= Delay1No60_out;
Delay1No61_out_to_Add22_impl_parent_implementedSystem_port_1_cast <= Delay1No61_out;
   Add22_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add22_impl_out,
                 X => Delay1No60_out_to_Add22_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No61_out_to_Add22_impl_parent_implementedSystem_port_1_cast);

SharedReg129_out_to_MUX_Add22_impl_0_parent_implementedSystem_port_1_cast <= SharedReg129_out;
SharedReg171_out_to_MUX_Add22_impl_0_parent_implementedSystem_port_2_cast <= SharedReg171_out;
   MUX_Add22_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg129_out_to_MUX_Add22_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg171_out_to_MUX_Add22_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add22_impl_0_out);

   Delay1No60_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add22_impl_0_out,
                 Y => Delay1No60_out);

SharedReg135_out_to_MUX_Add22_impl_1_parent_implementedSystem_port_1_cast <= SharedReg135_out;
SharedReg177_out_to_MUX_Add22_impl_1_parent_implementedSystem_port_2_cast <= SharedReg177_out;
   MUX_Add22_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg135_out_to_MUX_Add22_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg177_out_to_MUX_Add22_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add22_impl_1_out);

   Delay1No61_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add22_impl_1_out,
                 Y => Delay1No61_out);

Delay1No62_out_to_Add112_impl_parent_implementedSystem_port_0_cast <= Delay1No62_out;
Delay1No63_out_to_Add112_impl_parent_implementedSystem_port_1_cast <= Delay1No63_out;
   Add112_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add112_impl_out,
                 X => Delay1No62_out_to_Add112_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No63_out_to_Add112_impl_parent_implementedSystem_port_1_cast);

SharedReg118_out_to_MUX_Add112_impl_0_parent_implementedSystem_port_1_cast <= SharedReg118_out;
SharedReg166_out_to_MUX_Add112_impl_0_parent_implementedSystem_port_2_cast <= SharedReg166_out;
   MUX_Add112_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg118_out_to_MUX_Add112_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg166_out_to_MUX_Add112_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add112_impl_0_out);

   Delay1No62_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add112_impl_0_out,
                 Y => Delay1No62_out);

SharedReg130_out_to_MUX_Add112_impl_1_parent_implementedSystem_port_1_cast <= SharedReg130_out;
SharedReg172_out_to_MUX_Add112_impl_1_parent_implementedSystem_port_2_cast <= SharedReg172_out;
   MUX_Add112_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg130_out_to_MUX_Add112_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg172_out_to_MUX_Add112_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add112_impl_1_out);

   Delay1No63_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add112_impl_1_out,
                 Y => Delay1No63_out);

Delay1No64_out_to_Add24_impl_parent_implementedSystem_port_0_cast <= Delay1No64_out;
Delay1No65_out_to_Add24_impl_parent_implementedSystem_port_1_cast <= Delay1No65_out;
   Add24_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add24_impl_out,
                 X => Delay1No64_out_to_Add24_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No65_out_to_Add24_impl_parent_implementedSystem_port_1_cast);

SharedReg141_out_to_MUX_Add24_impl_0_parent_implementedSystem_port_1_cast <= SharedReg141_out;
SharedReg129_out_to_MUX_Add24_impl_0_parent_implementedSystem_port_2_cast <= SharedReg129_out;
   MUX_Add24_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg141_out_to_MUX_Add24_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg129_out_to_MUX_Add24_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add24_impl_0_out);

   Delay1No64_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add24_impl_0_out,
                 Y => Delay1No64_out);

SharedReg147_out_to_MUX_Add24_impl_1_parent_implementedSystem_port_1_cast <= SharedReg147_out;
SharedReg141_out_to_MUX_Add24_impl_1_parent_implementedSystem_port_2_cast <= SharedReg141_out;
   MUX_Add24_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg147_out_to_MUX_Add24_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg141_out_to_MUX_Add24_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add24_impl_1_out);

   Delay1No65_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add24_impl_1_out,
                 Y => Delay1No65_out);

Delay1No66_out_to_Add114_impl_parent_implementedSystem_port_0_cast <= Delay1No66_out;
Delay1No67_out_to_Add114_impl_parent_implementedSystem_port_1_cast <= Delay1No67_out;
   Add114_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add114_impl_out,
                 X => Delay1No66_out_to_Add114_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No67_out_to_Add114_impl_parent_implementedSystem_port_1_cast);

SharedReg136_out_to_MUX_Add114_impl_0_parent_implementedSystem_port_1_cast <= SharedReg136_out;
SharedReg124_out_to_MUX_Add114_impl_0_parent_implementedSystem_port_2_cast <= SharedReg124_out;
   MUX_Add114_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg136_out_to_MUX_Add114_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg124_out_to_MUX_Add114_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add114_impl_0_out);

   Delay1No66_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add114_impl_0_out,
                 Y => Delay1No66_out);

SharedReg142_out_to_MUX_Add114_impl_1_parent_implementedSystem_port_1_cast <= SharedReg142_out;
SharedReg136_out_to_MUX_Add114_impl_1_parent_implementedSystem_port_2_cast <= SharedReg136_out;
   MUX_Add114_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg142_out_to_MUX_Add114_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg136_out_to_MUX_Add114_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add114_impl_1_out);

   Delay1No67_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add114_impl_1_out,
                 Y => Delay1No67_out);

Delay1No68_out_to_Add25_impl_parent_implementedSystem_port_0_cast <= Delay1No68_out;
Delay1No69_out_to_Add25_impl_parent_implementedSystem_port_1_cast <= Delay1No69_out;
   Add25_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add25_impl_out,
                 X => Delay1No68_out_to_Add25_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No69_out_to_Add25_impl_parent_implementedSystem_port_1_cast);

SharedReg153_out_to_MUX_Add25_impl_0_parent_implementedSystem_port_1_cast <= SharedReg153_out;
SharedReg135_out_to_MUX_Add25_impl_0_parent_implementedSystem_port_2_cast <= SharedReg135_out;
   MUX_Add25_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg153_out_to_MUX_Add25_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg135_out_to_MUX_Add25_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add25_impl_0_out);

   Delay1No68_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add25_impl_0_out,
                 Y => Delay1No68_out);

SharedReg159_out_to_MUX_Add25_impl_1_parent_implementedSystem_port_1_cast <= SharedReg159_out;
SharedReg147_out_to_MUX_Add25_impl_1_parent_implementedSystem_port_2_cast <= SharedReg147_out;
   MUX_Add25_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg159_out_to_MUX_Add25_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg147_out_to_MUX_Add25_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add25_impl_1_out);

   Delay1No69_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add25_impl_1_out,
                 Y => Delay1No69_out);

Delay1No70_out_to_Add115_impl_parent_implementedSystem_port_0_cast <= Delay1No70_out;
Delay1No71_out_to_Add115_impl_parent_implementedSystem_port_1_cast <= Delay1No71_out;
   Add115_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add115_impl_out,
                 X => Delay1No70_out_to_Add115_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No71_out_to_Add115_impl_parent_implementedSystem_port_1_cast);

SharedReg148_out_to_MUX_Add115_impl_0_parent_implementedSystem_port_1_cast <= SharedReg148_out;
SharedReg130_out_to_MUX_Add115_impl_0_parent_implementedSystem_port_2_cast <= SharedReg130_out;
   MUX_Add115_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg148_out_to_MUX_Add115_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Add115_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add115_impl_0_out);

   Delay1No70_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add115_impl_0_out,
                 Y => Delay1No70_out);

SharedReg154_out_to_MUX_Add115_impl_1_parent_implementedSystem_port_1_cast <= SharedReg154_out;
SharedReg142_out_to_MUX_Add115_impl_1_parent_implementedSystem_port_2_cast <= SharedReg142_out;
   MUX_Add115_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg154_out_to_MUX_Add115_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg142_out_to_MUX_Add115_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add115_impl_1_out);

   Delay1No71_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add115_impl_1_out,
                 Y => Delay1No71_out);

Delay1No72_out_to_Add26_impl_parent_implementedSystem_port_0_cast <= Delay1No72_out;
Delay1No73_out_to_Add26_impl_parent_implementedSystem_port_1_cast <= Delay1No73_out;
   Add26_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add26_impl_out,
                 X => Delay1No72_out_to_Add26_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No73_out_to_Add26_impl_parent_implementedSystem_port_1_cast);

SharedReg183_out_to_MUX_Add26_impl_0_parent_implementedSystem_port_1_cast <= SharedReg183_out;
SharedReg153_out_to_MUX_Add26_impl_0_parent_implementedSystem_port_2_cast <= SharedReg153_out;
   MUX_Add26_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg183_out_to_MUX_Add26_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg153_out_to_MUX_Add26_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add26_impl_0_out);

   Delay1No72_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add26_impl_0_out,
                 Y => Delay1No72_out);

SharedReg189_out_to_MUX_Add26_impl_1_parent_implementedSystem_port_1_cast <= SharedReg189_out;
SharedReg189_out_to_MUX_Add26_impl_1_parent_implementedSystem_port_2_cast <= SharedReg189_out;
   MUX_Add26_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg189_out_to_MUX_Add26_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg189_out_to_MUX_Add26_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add26_impl_1_out);

   Delay1No73_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add26_impl_1_out,
                 Y => Delay1No73_out);

Delay1No74_out_to_Add116_impl_parent_implementedSystem_port_0_cast <= Delay1No74_out;
Delay1No75_out_to_Add116_impl_parent_implementedSystem_port_1_cast <= Delay1No75_out;
   Add116_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add116_impl_out,
                 X => Delay1No74_out_to_Add116_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No75_out_to_Add116_impl_parent_implementedSystem_port_1_cast);

SharedReg178_out_to_MUX_Add116_impl_0_parent_implementedSystem_port_1_cast <= SharedReg178_out;
SharedReg148_out_to_MUX_Add116_impl_0_parent_implementedSystem_port_2_cast <= SharedReg148_out;
   MUX_Add116_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg178_out_to_MUX_Add116_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg148_out_to_MUX_Add116_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add116_impl_0_out);

   Delay1No74_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add116_impl_0_out,
                 Y => Delay1No74_out);

SharedReg184_out_to_MUX_Add116_impl_1_parent_implementedSystem_port_1_cast <= SharedReg184_out;
SharedReg184_out_to_MUX_Add116_impl_1_parent_implementedSystem_port_2_cast <= SharedReg184_out;
   MUX_Add116_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg184_out_to_MUX_Add116_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg184_out_to_MUX_Add116_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add116_impl_1_out);

   Delay1No75_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add116_impl_1_out,
                 Y => Delay1No75_out);

Delay1No76_out_to_Add27_impl_parent_implementedSystem_port_0_cast <= Delay1No76_out;
Delay1No77_out_to_Add27_impl_parent_implementedSystem_port_1_cast <= Delay1No77_out;
   Add27_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add27_impl_out,
                 X => Delay1No76_out_to_Add27_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No77_out_to_Add27_impl_parent_implementedSystem_port_1_cast);

Delay2No6_out_to_MUX_Add27_impl_0_parent_implementedSystem_port_1_cast <= Delay2No6_out;
SharedReg159_out_to_MUX_Add27_impl_0_parent_implementedSystem_port_2_cast <= SharedReg159_out;
   MUX_Add27_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No6_out_to_MUX_Add27_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg159_out_to_MUX_Add27_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add27_impl_0_out);

   Delay1No76_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add27_impl_0_out,
                 Y => Delay1No76_out);

Delay2No14_out_to_MUX_Add27_impl_1_parent_implementedSystem_port_1_cast <= Delay2No14_out;
SharedReg195_out_to_MUX_Add27_impl_1_parent_implementedSystem_port_2_cast <= SharedReg195_out;
   MUX_Add27_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No14_out_to_MUX_Add27_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg195_out_to_MUX_Add27_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add27_impl_1_out);

   Delay1No77_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add27_impl_1_out,
                 Y => Delay1No77_out);

Delay1No78_out_to_Add117_impl_parent_implementedSystem_port_0_cast <= Delay1No78_out;
Delay1No79_out_to_Add117_impl_parent_implementedSystem_port_1_cast <= Delay1No79_out;
   Add117_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add117_impl_out,
                 X => Delay1No78_out_to_Add117_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No79_out_to_Add117_impl_parent_implementedSystem_port_1_cast);

SharedReg195_out_to_MUX_Add117_impl_0_parent_implementedSystem_port_1_cast <= SharedReg195_out;
SharedReg154_out_to_MUX_Add117_impl_0_parent_implementedSystem_port_2_cast <= SharedReg154_out;
   MUX_Add117_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg195_out_to_MUX_Add117_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg154_out_to_MUX_Add117_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add117_impl_0_out);

   Delay1No78_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add117_impl_0_out,
                 Y => Delay1No78_out);

SharedReg201_out_to_MUX_Add117_impl_1_parent_implementedSystem_port_1_cast <= SharedReg201_out;
SharedReg190_out_to_MUX_Add117_impl_1_parent_implementedSystem_port_2_cast <= SharedReg190_out;
   MUX_Add117_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg201_out_to_MUX_Add117_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg190_out_to_MUX_Add117_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add117_impl_1_out);

   Delay1No79_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add117_impl_1_out,
                 Y => Delay1No79_out);

Delay1No80_out_to_Add34_impl_parent_implementedSystem_port_0_cast <= Delay1No80_out;
Delay1No81_out_to_Add34_impl_parent_implementedSystem_port_1_cast <= Delay1No81_out;
   Add34_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add34_impl_out,
                 X => Delay1No80_out_to_Add34_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No81_out_to_Add34_impl_parent_implementedSystem_port_1_cast);

SharedReg190_out_to_MUX_Add34_impl_0_parent_implementedSystem_port_1_cast <= SharedReg190_out;
SharedReg6_out_to_MUX_Add34_impl_0_parent_implementedSystem_port_2_cast <= SharedReg6_out;
   MUX_Add34_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg190_out_to_MUX_Add34_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg6_out_to_MUX_Add34_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add34_impl_0_out);

   Delay1No80_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add34_impl_0_out,
                 Y => Delay1No80_out);

SharedReg196_out_to_MUX_Add34_impl_1_parent_implementedSystem_port_1_cast <= SharedReg196_out;
SharedReg22_out_to_MUX_Add34_impl_1_parent_implementedSystem_port_2_cast <= SharedReg22_out;
   MUX_Add34_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg196_out_to_MUX_Add34_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg22_out_to_MUX_Add34_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add34_impl_1_out);

   Delay1No81_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add34_impl_1_out,
                 Y => Delay1No81_out);

Delay1No82_out_to_Add124_impl_parent_implementedSystem_port_0_cast <= Delay1No82_out;
Delay1No83_out_to_Add124_impl_parent_implementedSystem_port_1_cast <= Delay1No83_out;
   Add124_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add124_impl_out,
                 X => Delay1No82_out_to_Add124_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No83_out_to_Add124_impl_parent_implementedSystem_port_1_cast);

SharedReg207_out_to_MUX_Add124_impl_0_parent_implementedSystem_port_1_cast <= SharedReg207_out;
SharedReg7_out_to_MUX_Add124_impl_0_parent_implementedSystem_port_2_cast <= SharedReg7_out;
   MUX_Add124_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg207_out_to_MUX_Add124_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg7_out_to_MUX_Add124_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add124_impl_0_out);

   Delay1No82_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add124_impl_0_out,
                 Y => Delay1No82_out);

SharedReg213_out_to_MUX_Add124_impl_1_parent_implementedSystem_port_1_cast <= SharedReg213_out;
SharedReg23_out_to_MUX_Add124_impl_1_parent_implementedSystem_port_2_cast <= SharedReg23_out;
   MUX_Add124_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg213_out_to_MUX_Add124_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg23_out_to_MUX_Add124_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add124_impl_1_out);

   Delay1No83_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add124_impl_1_out,
                 Y => Delay1No83_out);

Delay1No84_out_to_Add126_impl_parent_implementedSystem_port_0_cast <= Delay1No84_out;
Delay1No85_out_to_Add126_impl_parent_implementedSystem_port_1_cast <= Delay1No85_out;
   Add126_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add126_impl_out,
                 X => Delay1No84_out_to_Add126_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No85_out_to_Add126_impl_parent_implementedSystem_port_1_cast);

SharedReg202_out_to_MUX_Add126_impl_0_parent_implementedSystem_port_1_cast <= SharedReg202_out;
SharedReg10_out_to_MUX_Add126_impl_0_parent_implementedSystem_port_2_cast <= SharedReg10_out;
   MUX_Add126_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg202_out_to_MUX_Add126_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg10_out_to_MUX_Add126_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add126_impl_0_out);

   Delay1No84_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add126_impl_0_out,
                 Y => Delay1No84_out);

SharedReg208_out_to_MUX_Add126_impl_1_parent_implementedSystem_port_1_cast <= SharedReg208_out;
SharedReg26_out_to_MUX_Add126_impl_1_parent_implementedSystem_port_2_cast <= SharedReg26_out;
   MUX_Add126_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg208_out_to_MUX_Add126_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg26_out_to_MUX_Add126_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add126_impl_1_out);

   Delay1No85_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add126_impl_1_out,
                 Y => Delay1No85_out);

Delay1No86_out_to_Add37_impl_parent_implementedSystem_port_0_cast <= Delay1No86_out;
Delay1No87_out_to_Add37_impl_parent_implementedSystem_port_1_cast <= Delay1No87_out;
   Add37_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add37_impl_out,
                 X => Delay1No86_out_to_Add37_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No87_out_to_Add37_impl_parent_implementedSystem_port_1_cast);

Delay2No4_out_to_MUX_Add37_impl_0_parent_implementedSystem_port_1_cast <= Delay2No4_out;
SharedReg11_out_to_MUX_Add37_impl_0_parent_implementedSystem_port_2_cast <= SharedReg11_out;
   MUX_Add37_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No4_out_to_MUX_Add37_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg11_out_to_MUX_Add37_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add37_impl_0_out);

   Delay1No86_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add37_impl_0_out,
                 Y => Delay1No86_out);

Delay2No12_out_to_MUX_Add37_impl_1_parent_implementedSystem_port_1_cast <= Delay2No12_out;
SharedReg27_out_to_MUX_Add37_impl_1_parent_implementedSystem_port_2_cast <= SharedReg27_out;
   MUX_Add37_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No12_out_to_MUX_Add37_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg27_out_to_MUX_Add37_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add37_impl_1_out);

   Delay1No87_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add37_impl_1_out,
                 Y => Delay1No87_out);

Delay1No88_out_to_Add127_impl_parent_implementedSystem_port_0_cast <= Delay1No88_out;
Delay1No89_out_to_Add127_impl_parent_implementedSystem_port_1_cast <= Delay1No89_out;
   Add127_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add127_impl_out,
                 X => Delay1No88_out_to_Add127_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No89_out_to_Add127_impl_parent_implementedSystem_port_1_cast);

Delay2No5_out_to_MUX_Add127_impl_0_parent_implementedSystem_port_1_cast <= Delay2No5_out;
SharedReg14_out_to_MUX_Add127_impl_0_parent_implementedSystem_port_2_cast <= SharedReg14_out;
   MUX_Add127_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No5_out_to_MUX_Add127_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg14_out_to_MUX_Add127_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add127_impl_0_out);

   Delay1No88_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add127_impl_0_out,
                 Y => Delay1No88_out);

Delay2No13_out_to_MUX_Add127_impl_1_parent_implementedSystem_port_1_cast <= Delay2No13_out;
SharedReg30_out_to_MUX_Add127_impl_1_parent_implementedSystem_port_2_cast <= SharedReg30_out;
   MUX_Add127_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No13_out_to_MUX_Add127_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg30_out_to_MUX_Add127_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add127_impl_1_out);

   Delay1No89_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add127_impl_1_out,
                 Y => Delay1No89_out);

Delay1No90_out_to_Add129_impl_parent_implementedSystem_port_0_cast <= Delay1No90_out;
Delay1No91_out_to_Add129_impl_parent_implementedSystem_port_1_cast <= Delay1No91_out;
   Add129_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add129_impl_out,
                 X => Delay1No90_out_to_Add129_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No91_out_to_Add129_impl_parent_implementedSystem_port_1_cast);

Delay2No7_out_to_MUX_Add129_impl_0_parent_implementedSystem_port_1_cast <= Delay2No7_out;
SharedReg15_out_to_MUX_Add129_impl_0_parent_implementedSystem_port_2_cast <= SharedReg15_out;
   MUX_Add129_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No7_out_to_MUX_Add129_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg15_out_to_MUX_Add129_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add129_impl_0_out);

   Delay1No90_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add129_impl_0_out,
                 Y => Delay1No90_out);

Delay2No15_out_to_MUX_Add129_impl_1_parent_implementedSystem_port_1_cast <= Delay2No15_out;
SharedReg31_out_to_MUX_Add129_impl_1_parent_implementedSystem_port_2_cast <= SharedReg31_out;
   MUX_Add129_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No15_out_to_MUX_Add129_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg31_out_to_MUX_Add129_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add129_impl_1_out);

   Delay1No91_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add129_impl_1_out,
                 Y => Delay1No91_out);

Delay1No92_out_to_Add41_impl_parent_implementedSystem_port_0_cast <= Delay1No92_out;
Delay1No93_out_to_Add41_impl_parent_implementedSystem_port_1_cast <= Delay1No93_out;
   Add41_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add41_impl_out,
                 X => Delay1No92_out_to_Add41_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No93_out_to_Add41_impl_parent_implementedSystem_port_1_cast);

SharedReg81_out_to_MUX_Add41_impl_0_parent_implementedSystem_port_1_cast <= SharedReg81_out;
SharedReg83_out_to_MUX_Add41_impl_0_parent_implementedSystem_port_2_cast <= SharedReg83_out;
   MUX_Add41_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg81_out_to_MUX_Add41_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg83_out_to_MUX_Add41_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add41_impl_0_out);

   Delay1No92_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add41_impl_0_out,
                 Y => Delay1No92_out);

SharedReg165_out_to_MUX_Add41_impl_1_parent_implementedSystem_port_1_cast <= SharedReg165_out;
SharedReg214_out_to_MUX_Add41_impl_1_parent_implementedSystem_port_2_cast <= SharedReg214_out;
   MUX_Add41_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg165_out_to_MUX_Add41_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg214_out_to_MUX_Add41_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add41_impl_1_out);

   Delay1No93_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add41_impl_1_out,
                 Y => Delay1No93_out);

Delay1No94_out_to_Add131_impl_parent_implementedSystem_port_0_cast <= Delay1No94_out;
Delay1No95_out_to_Add131_impl_parent_implementedSystem_port_1_cast <= Delay1No95_out;
   Add131_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add131_impl_out,
                 X => Delay1No94_out_to_Add131_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No95_out_to_Add131_impl_parent_implementedSystem_port_1_cast);

SharedReg76_out_to_MUX_Add131_impl_0_parent_implementedSystem_port_1_cast <= SharedReg76_out;
SharedReg76_out_to_MUX_Add131_impl_0_parent_implementedSystem_port_2_cast <= SharedReg76_out;
   MUX_Add131_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg76_out_to_MUX_Add131_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg76_out_to_MUX_Add131_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add131_impl_0_out);

   Delay1No94_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add131_impl_0_out,
                 Y => Delay1No94_out);

SharedReg160_out_to_MUX_Add131_impl_1_parent_implementedSystem_port_1_cast <= SharedReg160_out;
SharedReg196_out_to_MUX_Add131_impl_1_parent_implementedSystem_port_2_cast <= SharedReg196_out;
   MUX_Add131_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg160_out_to_MUX_Add131_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg196_out_to_MUX_Add131_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add131_impl_1_out);

   Delay1No95_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add131_impl_1_out,
                 Y => Delay1No95_out);

Delay1No96_out_to_Add43_impl_parent_implementedSystem_port_0_cast <= Delay1No96_out;
Delay1No97_out_to_Add43_impl_parent_implementedSystem_port_1_cast <= Delay1No97_out;
   Add43_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add43_impl_out,
                 X => Delay1No96_out_to_Add43_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No97_out_to_Add43_impl_parent_implementedSystem_port_1_cast);

SharedReg79_out_to_MUX_Add43_impl_0_parent_implementedSystem_port_1_cast <= SharedReg79_out;
SharedReg78_out_to_MUX_Add43_impl_0_parent_implementedSystem_port_2_cast <= SharedReg78_out;
   MUX_Add43_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg79_out_to_MUX_Add43_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg78_out_to_MUX_Add43_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add43_impl_0_out);

   Delay1No96_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add43_impl_0_out,
                 Y => Delay1No96_out);

SharedReg80_out_to_MUX_Add43_impl_1_parent_implementedSystem_port_1_cast <= SharedReg80_out;
SharedReg79_out_to_MUX_Add43_impl_1_parent_implementedSystem_port_2_cast <= SharedReg79_out;
   MUX_Add43_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg80_out_to_MUX_Add43_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg79_out_to_MUX_Add43_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add43_impl_1_out);

   Delay1No97_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add43_impl_1_out,
                 Y => Delay1No97_out);

Delay1No98_out_to_Product4_impl_parent_implementedSystem_port_0_cast <= Delay1No98_out;
Delay1No99_out_to_Product4_impl_parent_implementedSystem_port_1_cast <= Delay1No99_out;
   Product4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_impl_out,
                 X => Delay1No98_out_to_Product4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No99_out_to_Product4_impl_parent_implementedSystem_port_1_cast);

SharedReg245_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg245_out;
SharedReg256_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg256_out;
   MUX_Product4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg245_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg256_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product4_impl_0_out);

   Delay1No98_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_impl_0_out,
                 Y => Delay1No98_out);

SharedReg263_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg263_out;
SharedReg32_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg32_out;
   MUX_Product4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg263_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg32_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product4_impl_1_out);

   Delay1No99_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_impl_1_out,
                 Y => Delay1No99_out);

Delay1No100_out_to_Product11_impl_parent_implementedSystem_port_0_cast <= Delay1No100_out;
Delay1No101_out_to_Product11_impl_parent_implementedSystem_port_1_cast <= Delay1No101_out;
   Product11_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product11_impl_out,
                 X => Delay1No100_out_to_Product11_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No101_out_to_Product11_impl_parent_implementedSystem_port_1_cast);

SharedReg258_out_to_MUX_Product11_impl_0_parent_implementedSystem_port_1_cast <= SharedReg258_out;
SharedReg256_out_to_MUX_Product11_impl_0_parent_implementedSystem_port_2_cast <= SharedReg256_out;
   MUX_Product11_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg258_out_to_MUX_Product11_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg256_out_to_MUX_Product11_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product11_impl_0_out);

   Delay1No100_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_impl_0_out,
                 Y => Delay1No100_out);

SharedReg33_out_to_MUX_Product11_impl_1_parent_implementedSystem_port_1_cast <= SharedReg33_out;
SharedReg33_out_to_MUX_Product11_impl_1_parent_implementedSystem_port_2_cast <= SharedReg33_out;
   MUX_Product11_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg33_out_to_MUX_Product11_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg33_out_to_MUX_Product11_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product11_impl_1_out);

   Delay1No101_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_impl_1_out,
                 Y => Delay1No101_out);

Delay1No102_out_to_Product21_impl_parent_implementedSystem_port_0_cast <= Delay1No102_out;
Delay1No103_out_to_Product21_impl_parent_implementedSystem_port_1_cast <= Delay1No103_out;
   Product21_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_impl_out,
                 X => Delay1No102_out_to_Product21_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No103_out_to_Product21_impl_parent_implementedSystem_port_1_cast);

SharedReg258_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_1_cast <= SharedReg258_out;
SharedReg257_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_2_cast <= SharedReg257_out;
   MUX_Product21_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg258_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg257_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product21_impl_0_out);

   Delay1No102_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_impl_0_out,
                 Y => Delay1No102_out);

SharedReg34_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_1_cast <= SharedReg34_out;
SharedReg32_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_2_cast <= SharedReg32_out;
   MUX_Product21_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg34_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg32_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product21_impl_1_out);

   Delay1No103_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_impl_1_out,
                 Y => Delay1No103_out);

Delay1No104_out_to_Product31_impl_parent_implementedSystem_port_0_cast <= Delay1No104_out;
Delay1No105_out_to_Product31_impl_parent_implementedSystem_port_1_cast <= Delay1No105_out;
   Product31_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product31_impl_out,
                 X => Delay1No104_out_to_Product31_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No105_out_to_Product31_impl_parent_implementedSystem_port_1_cast);

SharedReg259_out_to_MUX_Product31_impl_0_parent_implementedSystem_port_1_cast <= SharedReg259_out;
SharedReg33_out_to_MUX_Product31_impl_0_parent_implementedSystem_port_2_cast <= SharedReg33_out;
   MUX_Product31_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg259_out_to_MUX_Product31_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg33_out_to_MUX_Product31_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product31_impl_0_out);

   Delay1No104_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_impl_0_out,
                 Y => Delay1No104_out);

SharedReg33_out_to_MUX_Product31_impl_1_parent_implementedSystem_port_1_cast <= SharedReg33_out;
SharedReg257_out_to_MUX_Product31_impl_1_parent_implementedSystem_port_2_cast <= SharedReg257_out;
   MUX_Product31_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg33_out_to_MUX_Product31_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg257_out_to_MUX_Product31_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product31_impl_1_out);

   Delay1No105_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_impl_1_out,
                 Y => Delay1No105_out);

Delay1No106_out_to_Subtract2_impl_parent_implementedSystem_port_0_cast <= Delay1No106_out;
Delay1No107_out_to_Subtract2_impl_parent_implementedSystem_port_1_cast <= Delay1No107_out;
   Subtract2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_impl_out,
                 X => Delay1No106_out_to_Subtract2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No107_out_to_Subtract2_impl_parent_implementedSystem_port_1_cast);

SharedReg91_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg91_out;
SharedReg77_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg77_out;
   MUX_Subtract2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg91_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg77_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract2_impl_0_out);

   Delay1No106_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_impl_0_out,
                 Y => Delay1No106_out);

SharedReg77_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg77_out;
SharedReg80_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg80_out;
   MUX_Subtract2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg77_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg80_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract2_impl_1_out);

   Delay1No107_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_impl_1_out,
                 Y => Delay1No107_out);

Delay1No108_out_to_Product32_impl_parent_implementedSystem_port_0_cast <= Delay1No108_out;
Delay1No109_out_to_Product32_impl_parent_implementedSystem_port_1_cast <= Delay1No109_out;
   Product32_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_impl_out,
                 X => Delay1No108_out_to_Product32_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No109_out_to_Product32_impl_parent_implementedSystem_port_1_cast);

SharedReg34_out_to_MUX_Product32_impl_0_parent_implementedSystem_port_1_cast <= SharedReg34_out;
SharedReg272_out_to_MUX_Product32_impl_0_parent_implementedSystem_port_2_cast <= SharedReg272_out;
   MUX_Product32_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg34_out_to_MUX_Product32_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg272_out_to_MUX_Product32_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product32_impl_0_out);

   Delay1No108_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_impl_0_out,
                 Y => Delay1No108_out);

SharedReg259_out_to_MUX_Product32_impl_1_parent_implementedSystem_port_1_cast <= SharedReg259_out;
SharedReg74_out_to_MUX_Product32_impl_1_parent_implementedSystem_port_2_cast <= SharedReg74_out;
   MUX_Product32_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg259_out_to_MUX_Product32_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg74_out_to_MUX_Product32_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product32_impl_1_out);

   Delay1No109_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_impl_1_out,
                 Y => Delay1No109_out);

Delay1No110_out_to_Subtract3_impl_parent_implementedSystem_port_0_cast <= Delay1No110_out;
Delay1No111_out_to_Subtract3_impl_parent_implementedSystem_port_1_cast <= Delay1No111_out;
   Subtract3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract3_impl_out,
                 X => Delay1No110_out_to_Subtract3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No111_out_to_Subtract3_impl_parent_implementedSystem_port_1_cast);

SharedReg78_out_to_MUX_Subtract3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg78_out;
SharedReg82_out_to_MUX_Subtract3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg82_out;
   MUX_Subtract3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg78_out_to_MUX_Subtract3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg82_out_to_MUX_Subtract3_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract3_impl_0_out);

   Delay1No110_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_impl_0_out,
                 Y => Delay1No110_out);

SharedReg82_out_to_MUX_Subtract3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg82_out;
SharedReg87_out_to_MUX_Subtract3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg87_out;
   MUX_Subtract3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg82_out_to_MUX_Subtract3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg87_out_to_MUX_Subtract3_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract3_impl_1_out);

   Delay1No111_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_impl_1_out,
                 Y => Delay1No111_out);

Delay1No112_out_to_Add45_impl_parent_implementedSystem_port_0_cast <= Delay1No112_out;
Delay1No113_out_to_Add45_impl_parent_implementedSystem_port_1_cast <= Delay1No113_out;
   Add45_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add45_impl_out,
                 X => Delay1No112_out_to_Add45_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No113_out_to_Add45_impl_parent_implementedSystem_port_1_cast);

SharedReg86_out_to_MUX_Add45_impl_0_parent_implementedSystem_port_1_cast <= SharedReg86_out;
SharedReg85_out_to_MUX_Add45_impl_0_parent_implementedSystem_port_2_cast <= SharedReg85_out;
   MUX_Add45_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg86_out_to_MUX_Add45_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg85_out_to_MUX_Add45_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add45_impl_0_out);

   Delay1No112_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add45_impl_0_out,
                 Y => Delay1No112_out);

SharedReg87_out_to_MUX_Add45_impl_1_parent_implementedSystem_port_1_cast <= SharedReg87_out;
SharedReg86_out_to_MUX_Add45_impl_1_parent_implementedSystem_port_2_cast <= SharedReg86_out;
   MUX_Add45_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg87_out_to_MUX_Add45_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg86_out_to_MUX_Add45_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add45_impl_1_out);

   Delay1No113_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add45_impl_1_out,
                 Y => Delay1No113_out);

Delay1No114_out_to_Product6_impl_parent_implementedSystem_port_0_cast <= Delay1No114_out;
Delay1No115_out_to_Product6_impl_parent_implementedSystem_port_1_cast <= Delay1No115_out;
   Product6_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product6_impl_out,
                 X => Delay1No114_out_to_Product6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No115_out_to_Product6_impl_parent_implementedSystem_port_1_cast);

SharedReg260_out_to_MUX_Product6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg260_out;
SharedReg272_out_to_MUX_Product6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg272_out;
   MUX_Product6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg260_out_to_MUX_Product6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg272_out_to_MUX_Product6_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product6_impl_0_out);

   Delay1No114_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_impl_0_out,
                 Y => Delay1No114_out);

SharedReg238_out_to_MUX_Product6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg238_out;
SharedReg75_out_to_MUX_Product6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg75_out;
   MUX_Product6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg238_out_to_MUX_Product6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg75_out_to_MUX_Product6_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product6_impl_1_out);

   Delay1No115_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_impl_1_out,
                 Y => Delay1No115_out);

Delay1No116_out_to_Product13_impl_parent_implementedSystem_port_0_cast <= Delay1No116_out;
Delay1No117_out_to_Product13_impl_parent_implementedSystem_port_1_cast <= Delay1No117_out;
   Product13_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product13_impl_out,
                 X => Delay1No116_out_to_Product13_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No117_out_to_Product13_impl_parent_implementedSystem_port_1_cast);

SharedReg260_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_1_cast <= SharedReg260_out;
SharedReg273_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_2_cast <= SharedReg273_out;
   MUX_Product13_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg260_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg273_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product13_impl_0_out);

   Delay1No116_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product13_impl_0_out,
                 Y => Delay1No116_out);

SharedReg239_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_1_cast <= SharedReg239_out;
SharedReg74_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_2_cast <= SharedReg74_out;
   MUX_Product13_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg239_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg74_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product13_impl_1_out);

   Delay1No117_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product13_impl_1_out,
                 Y => Delay1No117_out);

Delay1No118_out_to_Product23_impl_parent_implementedSystem_port_0_cast <= Delay1No118_out;
Delay1No119_out_to_Product23_impl_parent_implementedSystem_port_1_cast <= Delay1No119_out;
   Product23_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product23_impl_out,
                 X => Delay1No118_out_to_Product23_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No119_out_to_Product23_impl_parent_implementedSystem_port_1_cast);

SharedReg261_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_1_cast <= SharedReg261_out;
SharedReg75_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_2_cast <= SharedReg75_out;
   MUX_Product23_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg261_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg75_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product23_impl_0_out);

   Delay1No118_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_impl_0_out,
                 Y => Delay1No118_out);

SharedReg238_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_1_cast <= SharedReg238_out;
SharedReg273_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_2_cast <= SharedReg273_out;
   MUX_Product23_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg238_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg273_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product23_impl_1_out);

   Delay1No119_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_impl_1_out,
                 Y => Delay1No119_out);

Delay1No120_out_to_Product33_impl_parent_implementedSystem_port_0_cast <= Delay1No120_out;
Delay1No121_out_to_Product33_impl_parent_implementedSystem_port_1_cast <= Delay1No121_out;
   Product33_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product33_impl_out,
                 X => Delay1No120_out_to_Product33_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No121_out_to_Product33_impl_parent_implementedSystem_port_1_cast);

SharedReg239_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_1_cast <= SharedReg239_out;
SharedReg291_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_2_cast <= SharedReg291_out;
   MUX_Product33_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg239_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg291_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product33_impl_0_out);

   Delay1No120_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_impl_0_out,
                 Y => Delay1No120_out);

SharedReg261_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_1_cast <= SharedReg261_out;
SharedReg34_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_2_cast <= SharedReg34_out;
   MUX_Product33_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg261_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg34_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product33_impl_1_out);

   Delay1No121_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_impl_1_out,
                 Y => Delay1No121_out);

Delay1No122_out_to_Subtract4_impl_parent_implementedSystem_port_0_cast <= Delay1No122_out;
Delay1No123_out_to_Subtract4_impl_parent_implementedSystem_port_1_cast <= Delay1No123_out;
   Subtract4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract4_impl_out,
                 X => Delay1No122_out_to_Subtract4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No123_out_to_Subtract4_impl_parent_implementedSystem_port_1_cast);

SharedReg85_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg85_out;
SharedReg92_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg92_out;
   MUX_Subtract4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg85_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg92_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract4_impl_0_out);

   Delay1No122_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_impl_0_out,
                 Y => Delay1No122_out);

SharedReg88_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg88_out;
SharedReg96_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg96_out;
   MUX_Subtract4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg88_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg96_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract4_impl_1_out);

   Delay1No123_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_impl_1_out,
                 Y => Delay1No123_out);

Delay1No124_out_to_Add46_impl_parent_implementedSystem_port_0_cast <= Delay1No124_out;
Delay1No125_out_to_Add46_impl_parent_implementedSystem_port_1_cast <= Delay1No125_out;
   Add46_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add46_impl_out,
                 X => Delay1No124_out_to_Add46_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No125_out_to_Add46_impl_parent_implementedSystem_port_1_cast);

SharedReg92_out_to_MUX_Add46_impl_0_parent_implementedSystem_port_1_cast <= SharedReg92_out;
SharedReg93_out_to_MUX_Add46_impl_0_parent_implementedSystem_port_2_cast <= SharedReg93_out;
   MUX_Add46_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg92_out_to_MUX_Add46_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg93_out_to_MUX_Add46_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add46_impl_0_out);

   Delay1No124_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add46_impl_0_out,
                 Y => Delay1No124_out);

SharedReg93_out_to_MUX_Add46_impl_1_parent_implementedSystem_port_1_cast <= SharedReg93_out;
SharedReg95_out_to_MUX_Add46_impl_1_parent_implementedSystem_port_2_cast <= SharedReg95_out;
   MUX_Add46_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg93_out_to_MUX_Add46_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg95_out_to_MUX_Add46_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add46_impl_1_out);

   Delay1No125_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add46_impl_1_out,
                 Y => Delay1No125_out);

Delay1No126_out_to_Product7_impl_parent_implementedSystem_port_0_cast <= Delay1No126_out;
Delay1No127_out_to_Product7_impl_parent_implementedSystem_port_1_cast <= Delay1No127_out;
   Product7_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product7_impl_out,
                 X => Delay1No126_out_to_Product7_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No127_out_to_Product7_impl_parent_implementedSystem_port_1_cast);

SharedReg262_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_1_cast <= SharedReg262_out;
SharedReg35_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_2_cast <= SharedReg35_out;
   MUX_Product7_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg262_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg35_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product7_impl_0_out);

   Delay1No126_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product7_impl_0_out,
                 Y => Delay1No126_out);

SharedReg244_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_1_cast <= SharedReg244_out;
SharedReg291_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_2_cast <= SharedReg291_out;
   MUX_Product7_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg244_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg291_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product7_impl_1_out);

   Delay1No127_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product7_impl_1_out,
                 Y => Delay1No127_out);

Delay1No128_out_to_Product14_impl_parent_implementedSystem_port_0_cast <= Delay1No128_out;
Delay1No129_out_to_Product14_impl_parent_implementedSystem_port_1_cast <= Delay1No129_out;
   Product14_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product14_impl_out,
                 X => Delay1No128_out_to_Product14_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No129_out_to_Product14_impl_parent_implementedSystem_port_1_cast);

SharedReg262_out_to_MUX_Product14_impl_0_parent_implementedSystem_port_1_cast <= SharedReg262_out;
SharedReg280_out_to_MUX_Product14_impl_0_parent_implementedSystem_port_2_cast <= SharedReg280_out;
   MUX_Product14_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg262_out_to_MUX_Product14_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg280_out_to_MUX_Product14_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product14_impl_0_out);

   Delay1No128_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product14_impl_0_out,
                 Y => Delay1No128_out);

SharedReg245_out_to_MUX_Product14_impl_1_parent_implementedSystem_port_1_cast <= SharedReg245_out;
SharedReg40_out_to_MUX_Product14_impl_1_parent_implementedSystem_port_2_cast <= SharedReg40_out;
   MUX_Product14_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg245_out_to_MUX_Product14_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg40_out_to_MUX_Product14_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product14_impl_1_out);

   Delay1No129_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product14_impl_1_out,
                 Y => Delay1No129_out);

Delay1No130_out_to_Product24_impl_parent_implementedSystem_port_0_cast <= Delay1No130_out;
Delay1No131_out_to_Product24_impl_parent_implementedSystem_port_1_cast <= Delay1No131_out;
   Product24_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product24_impl_out,
                 X => Delay1No130_out_to_Product24_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No131_out_to_Product24_impl_parent_implementedSystem_port_1_cast);

SharedReg263_out_to_MUX_Product24_impl_0_parent_implementedSystem_port_1_cast <= SharedReg263_out;
SharedReg280_out_to_MUX_Product24_impl_0_parent_implementedSystem_port_2_cast <= SharedReg280_out;
   MUX_Product24_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg263_out_to_MUX_Product24_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg280_out_to_MUX_Product24_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product24_impl_0_out);

   Delay1No130_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product24_impl_0_out,
                 Y => Delay1No130_out);

SharedReg244_out_to_MUX_Product24_impl_1_parent_implementedSystem_port_1_cast <= SharedReg244_out;
SharedReg41_out_to_MUX_Product24_impl_1_parent_implementedSystem_port_2_cast <= SharedReg41_out;
   MUX_Product24_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg244_out_to_MUX_Product24_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg41_out_to_MUX_Product24_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product24_impl_1_out);

   Delay1No131_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product24_impl_1_out,
                 Y => Delay1No131_out);

Delay1No132_out_to_Add47_impl_parent_implementedSystem_port_0_cast <= Delay1No132_out;
Delay1No133_out_to_Add47_impl_parent_implementedSystem_port_1_cast <= Delay1No133_out;
   Add47_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add47_impl_out,
                 X => Delay1No132_out_to_Add47_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No133_out_to_Add47_impl_parent_implementedSystem_port_1_cast);

SharedReg96_out_to_MUX_Add47_impl_0_parent_implementedSystem_port_1_cast <= SharedReg96_out;
SharedReg107_out_to_MUX_Add47_impl_0_parent_implementedSystem_port_2_cast <= SharedReg107_out;
   MUX_Add47_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg96_out_to_MUX_Add47_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg107_out_to_MUX_Add47_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add47_impl_0_out);

   Delay1No132_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add47_impl_0_out,
                 Y => Delay1No132_out);

SharedReg97_out_to_MUX_Add47_impl_1_parent_implementedSystem_port_1_cast <= SharedReg97_out;
SharedReg108_out_to_MUX_Add47_impl_1_parent_implementedSystem_port_2_cast <= SharedReg108_out;
   MUX_Add47_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg97_out_to_MUX_Add47_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg108_out_to_MUX_Add47_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add47_impl_1_out);

   Delay1No133_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add47_impl_1_out,
                 Y => Delay1No133_out);

Delay1No134_out_to_Product8_impl_parent_implementedSystem_port_0_cast <= Delay1No134_out;
Delay1No135_out_to_Product8_impl_parent_implementedSystem_port_1_cast <= Delay1No135_out;
   Product8_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product8_impl_out,
                 X => Delay1No134_out_to_Product8_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No135_out_to_Product8_impl_parent_implementedSystem_port_1_cast);

SharedReg264_out_to_MUX_Product8_impl_0_parent_implementedSystem_port_1_cast <= SharedReg264_out;
SharedReg281_out_to_MUX_Product8_impl_0_parent_implementedSystem_port_2_cast <= SharedReg281_out;
   MUX_Product8_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg264_out_to_MUX_Product8_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg281_out_to_MUX_Product8_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product8_impl_0_out);

   Delay1No134_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product8_impl_0_out,
                 Y => Delay1No134_out);

SharedReg246_out_to_MUX_Product8_impl_1_parent_implementedSystem_port_1_cast <= SharedReg246_out;
SharedReg40_out_to_MUX_Product8_impl_1_parent_implementedSystem_port_2_cast <= SharedReg40_out;
   MUX_Product8_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg246_out_to_MUX_Product8_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg40_out_to_MUX_Product8_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product8_impl_1_out);

   Delay1No135_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product8_impl_1_out,
                 Y => Delay1No135_out);

Delay1No136_out_to_Product15_impl_parent_implementedSystem_port_0_cast <= Delay1No136_out;
Delay1No137_out_to_Product15_impl_parent_implementedSystem_port_1_cast <= Delay1No137_out;
   Product15_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product15_impl_out,
                 X => Delay1No136_out_to_Product15_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No137_out_to_Product15_impl_parent_implementedSystem_port_1_cast);

SharedReg264_out_to_MUX_Product15_impl_0_parent_implementedSystem_port_1_cast <= SharedReg264_out;
SharedReg41_out_to_MUX_Product15_impl_0_parent_implementedSystem_port_2_cast <= SharedReg41_out;
   MUX_Product15_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg264_out_to_MUX_Product15_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg41_out_to_MUX_Product15_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product15_impl_0_out);

   Delay1No136_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product15_impl_0_out,
                 Y => Delay1No136_out);

SharedReg247_out_to_MUX_Product15_impl_1_parent_implementedSystem_port_1_cast <= SharedReg247_out;
SharedReg281_out_to_MUX_Product15_impl_1_parent_implementedSystem_port_2_cast <= SharedReg281_out;
   MUX_Product15_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg247_out_to_MUX_Product15_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg281_out_to_MUX_Product15_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product15_impl_1_out);

   Delay1No137_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product15_impl_1_out,
                 Y => Delay1No137_out);

Delay1No138_out_to_Product25_impl_parent_implementedSystem_port_0_cast <= Delay1No138_out;
Delay1No139_out_to_Product25_impl_parent_implementedSystem_port_1_cast <= Delay1No139_out;
   Product25_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product25_impl_out,
                 X => Delay1No138_out_to_Product25_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No139_out_to_Product25_impl_parent_implementedSystem_port_1_cast);

SharedReg265_out_to_MUX_Product25_impl_0_parent_implementedSystem_port_1_cast <= SharedReg265_out;
SharedReg290_out_to_MUX_Product25_impl_0_parent_implementedSystem_port_2_cast <= SharedReg290_out;
   MUX_Product25_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg265_out_to_MUX_Product25_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg290_out_to_MUX_Product25_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product25_impl_0_out);

   Delay1No138_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product25_impl_0_out,
                 Y => Delay1No138_out);

SharedReg246_out_to_MUX_Product25_impl_1_parent_implementedSystem_port_1_cast <= SharedReg246_out;
SharedReg34_out_to_MUX_Product25_impl_1_parent_implementedSystem_port_2_cast <= SharedReg34_out;
   MUX_Product25_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg246_out_to_MUX_Product25_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg34_out_to_MUX_Product25_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product25_impl_1_out);

   Delay1No139_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product25_impl_1_out,
                 Y => Delay1No139_out);

Delay1No140_out_to_Product35_impl_parent_implementedSystem_port_0_cast <= Delay1No140_out;
Delay1No141_out_to_Product35_impl_parent_implementedSystem_port_1_cast <= Delay1No141_out;
   Product35_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product35_impl_out,
                 X => Delay1No140_out_to_Product35_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No141_out_to_Product35_impl_parent_implementedSystem_port_1_cast);

SharedReg247_out_to_MUX_Product35_impl_0_parent_implementedSystem_port_1_cast <= SharedReg247_out;
SharedReg290_out_to_MUX_Product35_impl_0_parent_implementedSystem_port_2_cast <= SharedReg290_out;
   MUX_Product35_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg247_out_to_MUX_Product35_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg290_out_to_MUX_Product35_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product35_impl_0_out);

   Delay1No140_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product35_impl_0_out,
                 Y => Delay1No140_out);

SharedReg265_out_to_MUX_Product35_impl_1_parent_implementedSystem_port_1_cast <= SharedReg265_out;
SharedReg35_out_to_MUX_Product35_impl_1_parent_implementedSystem_port_2_cast <= SharedReg35_out;
   MUX_Product35_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg265_out_to_MUX_Product35_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg35_out_to_MUX_Product35_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product35_impl_1_out);

   Delay1No141_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product35_impl_1_out,
                 Y => Delay1No141_out);

Delay1No142_out_to_Subtract6_impl_parent_implementedSystem_port_0_cast <= Delay1No142_out;
Delay1No143_out_to_Subtract6_impl_parent_implementedSystem_port_1_cast <= Delay1No143_out;
   Subtract6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract6_impl_out,
                 X => Delay1No142_out_to_Subtract6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No143_out_to_Subtract6_impl_parent_implementedSystem_port_1_cast);

SharedReg95_out_to_MUX_Subtract6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg95_out;
SharedReg104_out_to_MUX_Subtract6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg104_out;
   MUX_Subtract6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg95_out_to_MUX_Subtract6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg104_out_to_MUX_Subtract6_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract6_impl_0_out);

   Delay1No142_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract6_impl_0_out,
                 Y => Delay1No142_out);

SharedReg98_out_to_MUX_Subtract6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg98_out;
SharedReg109_out_to_MUX_Subtract6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg109_out;
   MUX_Subtract6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg98_out_to_MUX_Subtract6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg109_out_to_MUX_Subtract6_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract6_impl_1_out);

   Delay1No143_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract6_impl_1_out,
                 Y => Delay1No143_out);

Delay1No144_out_to_Add48_impl_parent_implementedSystem_port_0_cast <= Delay1No144_out;
Delay1No145_out_to_Add48_impl_parent_implementedSystem_port_1_cast <= Delay1No145_out;
   Add48_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add48_impl_out,
                 X => Delay1No144_out_to_Add48_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No145_out_to_Add48_impl_parent_implementedSystem_port_1_cast);

SharedReg102_out_to_MUX_Add48_impl_0_parent_implementedSystem_port_1_cast <= SharedReg102_out;
SharedReg113_out_to_MUX_Add48_impl_0_parent_implementedSystem_port_2_cast <= SharedReg113_out;
   MUX_Add48_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg102_out_to_MUX_Add48_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg113_out_to_MUX_Add48_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add48_impl_0_out);

   Delay1No144_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add48_impl_0_out,
                 Y => Delay1No144_out);

SharedReg103_out_to_MUX_Add48_impl_1_parent_implementedSystem_port_1_cast <= SharedReg103_out;
SharedReg114_out_to_MUX_Add48_impl_1_parent_implementedSystem_port_2_cast <= SharedReg114_out;
   MUX_Add48_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg103_out_to_MUX_Add48_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg114_out_to_MUX_Add48_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add48_impl_1_out);

   Delay1No145_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add48_impl_1_out,
                 Y => Delay1No145_out);

Delay1No146_out_to_Product9_impl_parent_implementedSystem_port_0_cast <= Delay1No146_out;
Delay1No147_out_to_Product9_impl_parent_implementedSystem_port_1_cast <= Delay1No147_out;
   Product9_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product9_impl_out,
                 X => Delay1No146_out_to_Product9_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No147_out_to_Product9_impl_parent_implementedSystem_port_1_cast);

SharedReg266_out_to_MUX_Product9_impl_0_parent_implementedSystem_port_1_cast <= SharedReg266_out;
SharedReg310_out_to_MUX_Product9_impl_0_parent_implementedSystem_port_2_cast <= SharedReg310_out;
   MUX_Product9_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg266_out_to_MUX_Product9_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg310_out_to_MUX_Product9_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product9_impl_0_out);

   Delay1No146_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product9_impl_0_out,
                 Y => Delay1No146_out);

SharedReg248_out_to_MUX_Product9_impl_1_parent_implementedSystem_port_1_cast <= SharedReg248_out;
SharedReg45_out_to_MUX_Product9_impl_1_parent_implementedSystem_port_2_cast <= SharedReg45_out;
   MUX_Product9_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg248_out_to_MUX_Product9_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg45_out_to_MUX_Product9_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product9_impl_1_out);

   Delay1No147_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product9_impl_1_out,
                 Y => Delay1No147_out);

Delay1No148_out_to_Product16_impl_parent_implementedSystem_port_0_cast <= Delay1No148_out;
Delay1No149_out_to_Product16_impl_parent_implementedSystem_port_1_cast <= Delay1No149_out;
   Product16_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product16_impl_out,
                 X => Delay1No148_out_to_Product16_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No149_out_to_Product16_impl_parent_implementedSystem_port_1_cast);

SharedReg266_out_to_MUX_Product16_impl_0_parent_implementedSystem_port_1_cast <= SharedReg266_out;
SharedReg310_out_to_MUX_Product16_impl_0_parent_implementedSystem_port_2_cast <= SharedReg310_out;
   MUX_Product16_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg266_out_to_MUX_Product16_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg310_out_to_MUX_Product16_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product16_impl_0_out);

   Delay1No148_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product16_impl_0_out,
                 Y => Delay1No148_out);

SharedReg249_out_to_MUX_Product16_impl_1_parent_implementedSystem_port_1_cast <= SharedReg249_out;
SharedReg47_out_to_MUX_Product16_impl_1_parent_implementedSystem_port_2_cast <= SharedReg47_out;
   MUX_Product16_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg249_out_to_MUX_Product16_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg47_out_to_MUX_Product16_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product16_impl_1_out);

   Delay1No149_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product16_impl_1_out,
                 Y => Delay1No149_out);

Delay1No150_out_to_Product26_impl_parent_implementedSystem_port_0_cast <= Delay1No150_out;
Delay1No151_out_to_Product26_impl_parent_implementedSystem_port_1_cast <= Delay1No151_out;
   Product26_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product26_impl_out,
                 X => Delay1No150_out_to_Product26_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No151_out_to_Product26_impl_parent_implementedSystem_port_1_cast);

SharedReg267_out_to_MUX_Product26_impl_0_parent_implementedSystem_port_1_cast <= SharedReg267_out;
SharedReg311_out_to_MUX_Product26_impl_0_parent_implementedSystem_port_2_cast <= SharedReg311_out;
   MUX_Product26_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg267_out_to_MUX_Product26_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg311_out_to_MUX_Product26_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product26_impl_0_out);

   Delay1No150_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product26_impl_0_out,
                 Y => Delay1No150_out);

SharedReg248_out_to_MUX_Product26_impl_1_parent_implementedSystem_port_1_cast <= SharedReg248_out;
SharedReg45_out_to_MUX_Product26_impl_1_parent_implementedSystem_port_2_cast <= SharedReg45_out;
   MUX_Product26_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg248_out_to_MUX_Product26_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg45_out_to_MUX_Product26_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product26_impl_1_out);

   Delay1No151_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product26_impl_1_out,
                 Y => Delay1No151_out);

Delay1No152_out_to_Product36_impl_parent_implementedSystem_port_0_cast <= Delay1No152_out;
Delay1No153_out_to_Product36_impl_parent_implementedSystem_port_1_cast <= Delay1No153_out;
   Product36_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product36_impl_out,
                 X => Delay1No152_out_to_Product36_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No153_out_to_Product36_impl_parent_implementedSystem_port_1_cast);

SharedReg249_out_to_MUX_Product36_impl_0_parent_implementedSystem_port_1_cast <= SharedReg249_out;
SharedReg294_out_to_MUX_Product36_impl_0_parent_implementedSystem_port_2_cast <= SharedReg294_out;
   MUX_Product36_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg249_out_to_MUX_Product36_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg294_out_to_MUX_Product36_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product36_impl_0_out);

   Delay1No152_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product36_impl_0_out,
                 Y => Delay1No152_out);

SharedReg267_out_to_MUX_Product36_impl_1_parent_implementedSystem_port_1_cast <= SharedReg267_out;
SharedReg254_out_to_MUX_Product36_impl_1_parent_implementedSystem_port_2_cast <= SharedReg254_out;
   MUX_Product36_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg267_out_to_MUX_Product36_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg254_out_to_MUX_Product36_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product36_impl_1_out);

   Delay1No153_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product36_impl_1_out,
                 Y => Delay1No153_out);

Delay1No154_out_to_Subtract7_impl_parent_implementedSystem_port_0_cast <= Delay1No154_out;
Delay1No155_out_to_Subtract7_impl_parent_implementedSystem_port_1_cast <= Delay1No155_out;
   Subtract7_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract7_impl_out,
                 X => Delay1No154_out_to_Subtract7_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No155_out_to_Subtract7_impl_parent_implementedSystem_port_1_cast);

SharedReg101_out_to_MUX_Subtract7_impl_0_parent_implementedSystem_port_1_cast <= SharedReg101_out;
SharedReg110_out_to_MUX_Subtract7_impl_0_parent_implementedSystem_port_2_cast <= SharedReg110_out;
   MUX_Subtract7_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg101_out_to_MUX_Subtract7_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg110_out_to_MUX_Subtract7_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract7_impl_0_out);

   Delay1No154_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract7_impl_0_out,
                 Y => Delay1No154_out);

SharedReg104_out_to_MUX_Subtract7_impl_1_parent_implementedSystem_port_1_cast <= SharedReg104_out;
SharedReg115_out_to_MUX_Subtract7_impl_1_parent_implementedSystem_port_2_cast <= SharedReg115_out;
   MUX_Subtract7_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg104_out_to_MUX_Subtract7_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg115_out_to_MUX_Subtract7_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract7_impl_1_out);

   Delay1No155_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract7_impl_1_out,
                 Y => Delay1No155_out);

Delay1No156_out_to_Add49_impl_parent_implementedSystem_port_0_cast <= Delay1No156_out;
Delay1No157_out_to_Add49_impl_parent_implementedSystem_port_1_cast <= Delay1No157_out;
   Add49_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add49_impl_out,
                 X => Delay1No156_out_to_Add49_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No157_out_to_Add49_impl_parent_implementedSystem_port_1_cast);

SharedReg108_out_to_MUX_Add49_impl_0_parent_implementedSystem_port_1_cast <= SharedReg108_out;
SharedReg119_out_to_MUX_Add49_impl_0_parent_implementedSystem_port_2_cast <= SharedReg119_out;
   MUX_Add49_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg108_out_to_MUX_Add49_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg119_out_to_MUX_Add49_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add49_impl_0_out);

   Delay1No156_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add49_impl_0_out,
                 Y => Delay1No156_out);

SharedReg109_out_to_MUX_Add49_impl_1_parent_implementedSystem_port_1_cast <= SharedReg109_out;
SharedReg120_out_to_MUX_Add49_impl_1_parent_implementedSystem_port_2_cast <= SharedReg120_out;
   MUX_Add49_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg109_out_to_MUX_Add49_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg120_out_to_MUX_Add49_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add49_impl_1_out);

   Delay1No157_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add49_impl_1_out,
                 Y => Delay1No157_out);

Delay1No158_out_to_Product10_impl_parent_implementedSystem_port_0_cast <= Delay1No158_out;
Delay1No159_out_to_Product10_impl_parent_implementedSystem_port_1_cast <= Delay1No159_out;
   Product10_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product10_impl_out,
                 X => Delay1No158_out_to_Product10_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No159_out_to_Product10_impl_parent_implementedSystem_port_1_cast);

SharedReg300_out_to_MUX_Product10_impl_0_parent_implementedSystem_port_1_cast <= SharedReg300_out;
SharedReg294_out_to_MUX_Product10_impl_0_parent_implementedSystem_port_2_cast <= SharedReg294_out;
   MUX_Product10_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg300_out_to_MUX_Product10_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg294_out_to_MUX_Product10_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product10_impl_0_out);

   Delay1No158_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product10_impl_0_out,
                 Y => Delay1No158_out);

SharedReg250_out_to_MUX_Product10_impl_1_parent_implementedSystem_port_1_cast <= SharedReg250_out;
SharedReg255_out_to_MUX_Product10_impl_1_parent_implementedSystem_port_2_cast <= SharedReg255_out;
   MUX_Product10_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg250_out_to_MUX_Product10_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg255_out_to_MUX_Product10_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product10_impl_1_out);

   Delay1No159_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product10_impl_1_out,
                 Y => Delay1No159_out);

Delay1No160_out_to_Product17_impl_parent_implementedSystem_port_0_cast <= Delay1No160_out;
Delay1No161_out_to_Product17_impl_parent_implementedSystem_port_1_cast <= Delay1No161_out;
   Product17_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product17_impl_out,
                 X => Delay1No160_out_to_Product17_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No161_out_to_Product17_impl_parent_implementedSystem_port_1_cast);

SharedReg300_out_to_MUX_Product17_impl_0_parent_implementedSystem_port_1_cast <= SharedReg300_out;
SharedReg295_out_to_MUX_Product17_impl_0_parent_implementedSystem_port_2_cast <= SharedReg295_out;
   MUX_Product17_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg300_out_to_MUX_Product17_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg295_out_to_MUX_Product17_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product17_impl_0_out);

   Delay1No160_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product17_impl_0_out,
                 Y => Delay1No160_out);

SharedReg251_out_to_MUX_Product17_impl_1_parent_implementedSystem_port_1_cast <= SharedReg251_out;
SharedReg254_out_to_MUX_Product17_impl_1_parent_implementedSystem_port_2_cast <= SharedReg254_out;
   MUX_Product17_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg251_out_to_MUX_Product17_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg254_out_to_MUX_Product17_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product17_impl_1_out);

   Delay1No161_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product17_impl_1_out,
                 Y => Delay1No161_out);

Delay1No162_out_to_Product27_impl_parent_implementedSystem_port_0_cast <= Delay1No162_out;
Delay1No163_out_to_Product27_impl_parent_implementedSystem_port_1_cast <= Delay1No163_out;
   Product27_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product27_impl_out,
                 X => Delay1No162_out_to_Product27_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No163_out_to_Product27_impl_parent_implementedSystem_port_1_cast);

SharedReg301_out_to_MUX_Product27_impl_0_parent_implementedSystem_port_1_cast <= SharedReg301_out;
SharedReg255_out_to_MUX_Product27_impl_0_parent_implementedSystem_port_2_cast <= SharedReg255_out;
   MUX_Product27_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg301_out_to_MUX_Product27_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg255_out_to_MUX_Product27_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product27_impl_0_out);

   Delay1No162_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product27_impl_0_out,
                 Y => Delay1No162_out);

SharedReg250_out_to_MUX_Product27_impl_1_parent_implementedSystem_port_1_cast <= SharedReg250_out;
SharedReg295_out_to_MUX_Product27_impl_1_parent_implementedSystem_port_2_cast <= SharedReg295_out;
   MUX_Product27_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg250_out_to_MUX_Product27_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg295_out_to_MUX_Product27_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product27_impl_1_out);

   Delay1No163_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product27_impl_1_out,
                 Y => Delay1No163_out);

Delay1No164_out_to_Product37_impl_parent_implementedSystem_port_0_cast <= Delay1No164_out;
Delay1No165_out_to_Product37_impl_parent_implementedSystem_port_1_cast <= Delay1No165_out;
   Product37_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product37_impl_out,
                 X => Delay1No164_out_to_Product37_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No165_out_to_Product37_impl_parent_implementedSystem_port_1_cast);

SharedReg251_out_to_MUX_Product37_impl_0_parent_implementedSystem_port_1_cast <= SharedReg251_out;
SharedReg306_out_to_MUX_Product37_impl_0_parent_implementedSystem_port_2_cast <= SharedReg306_out;
   MUX_Product37_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg251_out_to_MUX_Product37_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg306_out_to_MUX_Product37_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product37_impl_0_out);

   Delay1No164_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product37_impl_0_out,
                 Y => Delay1No164_out);

SharedReg301_out_to_MUX_Product37_impl_1_parent_implementedSystem_port_1_cast <= SharedReg301_out;
SharedReg225_out_to_MUX_Product37_impl_1_parent_implementedSystem_port_2_cast <= SharedReg225_out;
   MUX_Product37_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg301_out_to_MUX_Product37_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg225_out_to_MUX_Product37_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product37_impl_1_out);

   Delay1No165_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product37_impl_1_out,
                 Y => Delay1No165_out);

Delay1No166_out_to_Subtract8_impl_parent_implementedSystem_port_0_cast <= Delay1No166_out;
Delay1No167_out_to_Subtract8_impl_parent_implementedSystem_port_1_cast <= Delay1No167_out;
   Subtract8_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract8_impl_out,
                 X => Delay1No166_out_to_Subtract8_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No167_out_to_Subtract8_impl_parent_implementedSystem_port_1_cast);

SharedReg107_out_to_MUX_Subtract8_impl_0_parent_implementedSystem_port_1_cast <= SharedReg107_out;
SharedReg116_out_to_MUX_Subtract8_impl_0_parent_implementedSystem_port_2_cast <= SharedReg116_out;
   MUX_Subtract8_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg107_out_to_MUX_Subtract8_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg116_out_to_MUX_Subtract8_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract8_impl_0_out);

   Delay1No166_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract8_impl_0_out,
                 Y => Delay1No166_out);

SharedReg110_out_to_MUX_Subtract8_impl_1_parent_implementedSystem_port_1_cast <= SharedReg110_out;
SharedReg121_out_to_MUX_Subtract8_impl_1_parent_implementedSystem_port_2_cast <= SharedReg121_out;
   MUX_Subtract8_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg110_out_to_MUX_Subtract8_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg121_out_to_MUX_Subtract8_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract8_impl_1_out);

   Delay1No167_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract8_impl_1_out,
                 Y => Delay1No167_out);

Delay1No168_out_to_Add50_impl_parent_implementedSystem_port_0_cast <= Delay1No168_out;
Delay1No169_out_to_Add50_impl_parent_implementedSystem_port_1_cast <= Delay1No169_out;
   Add50_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add50_impl_out,
                 X => Delay1No168_out_to_Add50_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No169_out_to_Add50_impl_parent_implementedSystem_port_1_cast);

SharedReg114_out_to_MUX_Add50_impl_0_parent_implementedSystem_port_1_cast <= SharedReg114_out;
SharedReg102_out_to_MUX_Add50_impl_0_parent_implementedSystem_port_2_cast <= SharedReg102_out;
   MUX_Add50_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg114_out_to_MUX_Add50_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg102_out_to_MUX_Add50_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add50_impl_0_out);

   Delay1No168_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add50_impl_0_out,
                 Y => Delay1No168_out);

SharedReg115_out_to_MUX_Add50_impl_1_parent_implementedSystem_port_1_cast <= SharedReg115_out;
SharedReg103_out_to_MUX_Add50_impl_1_parent_implementedSystem_port_2_cast <= SharedReg103_out;
   MUX_Add50_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg115_out_to_MUX_Add50_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg103_out_to_MUX_Add50_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add50_impl_1_out);

   Delay1No169_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add50_impl_1_out,
                 Y => Delay1No169_out);

Delay1No170_out_to_Product18_impl_parent_implementedSystem_port_0_cast <= Delay1No170_out;
Delay1No171_out_to_Product18_impl_parent_implementedSystem_port_1_cast <= Delay1No171_out;
   Product18_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product18_impl_out,
                 X => Delay1No170_out_to_Product18_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No171_out_to_Product18_impl_parent_implementedSystem_port_1_cast);

SharedReg270_out_to_MUX_Product18_impl_0_parent_implementedSystem_port_1_cast <= SharedReg270_out;
SharedReg306_out_to_MUX_Product18_impl_0_parent_implementedSystem_port_2_cast <= SharedReg306_out;
   MUX_Product18_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg270_out_to_MUX_Product18_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg306_out_to_MUX_Product18_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product18_impl_0_out);

   Delay1No170_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product18_impl_0_out,
                 Y => Delay1No170_out);

SharedReg252_out_to_MUX_Product18_impl_1_parent_implementedSystem_port_1_cast <= SharedReg252_out;
SharedReg226_out_to_MUX_Product18_impl_1_parent_implementedSystem_port_2_cast <= SharedReg226_out;
   MUX_Product18_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg252_out_to_MUX_Product18_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg226_out_to_MUX_Product18_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product18_impl_1_out);

   Delay1No171_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product18_impl_1_out,
                 Y => Delay1No171_out);

Delay1No172_out_to_Product19_impl_parent_implementedSystem_port_0_cast <= Delay1No172_out;
Delay1No173_out_to_Product19_impl_parent_implementedSystem_port_1_cast <= Delay1No173_out;
   Product19_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product19_impl_out,
                 X => Delay1No172_out_to_Product19_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No173_out_to_Product19_impl_parent_implementedSystem_port_1_cast);

SharedReg270_out_to_MUX_Product19_impl_0_parent_implementedSystem_port_1_cast <= SharedReg270_out;
SharedReg307_out_to_MUX_Product19_impl_0_parent_implementedSystem_port_2_cast <= SharedReg307_out;
   MUX_Product19_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg270_out_to_MUX_Product19_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg307_out_to_MUX_Product19_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product19_impl_0_out);

   Delay1No172_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product19_impl_0_out,
                 Y => Delay1No172_out);

SharedReg253_out_to_MUX_Product19_impl_1_parent_implementedSystem_port_1_cast <= SharedReg253_out;
SharedReg225_out_to_MUX_Product19_impl_1_parent_implementedSystem_port_2_cast <= SharedReg225_out;
   MUX_Product19_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg253_out_to_MUX_Product19_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg225_out_to_MUX_Product19_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product19_impl_1_out);

   Delay1No173_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product19_impl_1_out,
                 Y => Delay1No173_out);

Delay1No174_out_to_Product28_impl_parent_implementedSystem_port_0_cast <= Delay1No174_out;
Delay1No175_out_to_Product28_impl_parent_implementedSystem_port_1_cast <= Delay1No175_out;
   Product28_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product28_impl_out,
                 X => Delay1No174_out_to_Product28_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No175_out_to_Product28_impl_parent_implementedSystem_port_1_cast);

SharedReg271_out_to_MUX_Product28_impl_0_parent_implementedSystem_port_1_cast <= SharedReg271_out;
SharedReg226_out_to_MUX_Product28_impl_0_parent_implementedSystem_port_2_cast <= SharedReg226_out;
   MUX_Product28_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg271_out_to_MUX_Product28_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg226_out_to_MUX_Product28_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product28_impl_0_out);

   Delay1No174_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_impl_0_out,
                 Y => Delay1No174_out);

SharedReg252_out_to_MUX_Product28_impl_1_parent_implementedSystem_port_1_cast <= SharedReg252_out;
SharedReg307_out_to_MUX_Product28_impl_1_parent_implementedSystem_port_2_cast <= SharedReg307_out;
   MUX_Product28_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg252_out_to_MUX_Product28_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg307_out_to_MUX_Product28_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product28_impl_1_out);

   Delay1No175_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_impl_1_out,
                 Y => Delay1No175_out);

Delay1No176_out_to_Product38_impl_parent_implementedSystem_port_0_cast <= Delay1No176_out;
Delay1No177_out_to_Product38_impl_parent_implementedSystem_port_1_cast <= Delay1No177_out;
   Product38_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product38_impl_out,
                 X => Delay1No176_out_to_Product38_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No177_out_to_Product38_impl_parent_implementedSystem_port_1_cast);

SharedReg253_out_to_MUX_Product38_impl_0_parent_implementedSystem_port_1_cast <= SharedReg253_out;
SharedReg308_out_to_MUX_Product38_impl_0_parent_implementedSystem_port_2_cast <= SharedReg308_out;
   MUX_Product38_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg253_out_to_MUX_Product38_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg308_out_to_MUX_Product38_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product38_impl_0_out);

   Delay1No176_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product38_impl_0_out,
                 Y => Delay1No176_out);

SharedReg271_out_to_MUX_Product38_impl_1_parent_implementedSystem_port_1_cast <= SharedReg271_out;
SharedReg36_out_to_MUX_Product38_impl_1_parent_implementedSystem_port_2_cast <= SharedReg36_out;
   MUX_Product38_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg271_out_to_MUX_Product38_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg36_out_to_MUX_Product38_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product38_impl_1_out);

   Delay1No177_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product38_impl_1_out,
                 Y => Delay1No177_out);

Delay1No178_out_to_Subtract9_impl_parent_implementedSystem_port_0_cast <= Delay1No178_out;
Delay1No179_out_to_Subtract9_impl_parent_implementedSystem_port_1_cast <= Delay1No179_out;
   Subtract9_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract9_impl_out,
                 X => Delay1No178_out_to_Subtract9_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No179_out_to_Subtract9_impl_parent_implementedSystem_port_1_cast);

SharedReg113_out_to_MUX_Subtract9_impl_0_parent_implementedSystem_port_1_cast <= SharedReg113_out;
SharedReg101_out_to_MUX_Subtract9_impl_0_parent_implementedSystem_port_2_cast <= SharedReg101_out;
   MUX_Subtract9_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg113_out_to_MUX_Subtract9_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg101_out_to_MUX_Subtract9_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract9_impl_0_out);

   Delay1No178_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_impl_0_out,
                 Y => Delay1No178_out);

SharedReg116_out_to_MUX_Subtract9_impl_1_parent_implementedSystem_port_1_cast <= SharedReg116_out;
SharedReg128_out_to_MUX_Subtract9_impl_1_parent_implementedSystem_port_2_cast <= SharedReg128_out;
   MUX_Subtract9_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg116_out_to_MUX_Subtract9_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg128_out_to_MUX_Subtract9_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract9_impl_1_out);

   Delay1No179_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_impl_1_out,
                 Y => Delay1No179_out);

Delay1No180_out_to_Add52_impl_parent_implementedSystem_port_0_cast <= Delay1No180_out;
Delay1No181_out_to_Add52_impl_parent_implementedSystem_port_1_cast <= Delay1No181_out;
   Add52_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add52_impl_out,
                 X => Delay1No180_out_to_Add52_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No181_out_to_Add52_impl_parent_implementedSystem_port_1_cast);

SharedReg120_out_to_MUX_Add52_impl_0_parent_implementedSystem_port_1_cast <= SharedReg120_out;
SharedReg132_out_to_MUX_Add52_impl_0_parent_implementedSystem_port_2_cast <= SharedReg132_out;
   MUX_Add52_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg120_out_to_MUX_Add52_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg132_out_to_MUX_Add52_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add52_impl_0_out);

   Delay1No180_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add52_impl_0_out,
                 Y => Delay1No180_out);

SharedReg121_out_to_MUX_Add52_impl_1_parent_implementedSystem_port_1_cast <= SharedReg121_out;
SharedReg133_out_to_MUX_Add52_impl_1_parent_implementedSystem_port_2_cast <= SharedReg133_out;
   MUX_Add52_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg121_out_to_MUX_Add52_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg133_out_to_MUX_Add52_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add52_impl_1_out);

   Delay1No181_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add52_impl_1_out,
                 Y => Delay1No181_out);

Delay1No182_out_to_Product30_impl_parent_implementedSystem_port_0_cast <= Delay1No182_out;
Delay1No183_out_to_Product30_impl_parent_implementedSystem_port_1_cast <= Delay1No183_out;
   Product30_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product30_impl_out,
                 X => Delay1No182_out_to_Product30_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No183_out_to_Product30_impl_parent_implementedSystem_port_1_cast);

SharedReg274_out_to_MUX_Product30_impl_0_parent_implementedSystem_port_1_cast <= SharedReg274_out;
SharedReg308_out_to_MUX_Product30_impl_0_parent_implementedSystem_port_2_cast <= SharedReg308_out;
   MUX_Product30_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg274_out_to_MUX_Product30_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg308_out_to_MUX_Product30_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product30_impl_0_out);

   Delay1No182_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product30_impl_0_out,
                 Y => Delay1No182_out);

SharedReg74_out_to_MUX_Product30_impl_1_parent_implementedSystem_port_1_cast <= SharedReg74_out;
SharedReg37_out_to_MUX_Product30_impl_1_parent_implementedSystem_port_2_cast <= SharedReg37_out;
   MUX_Product30_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg74_out_to_MUX_Product30_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg37_out_to_MUX_Product30_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product30_impl_1_out);

   Delay1No183_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product30_impl_1_out,
                 Y => Delay1No183_out);

Delay1No184_out_to_Product111_impl_parent_implementedSystem_port_0_cast <= Delay1No184_out;
Delay1No185_out_to_Product111_impl_parent_implementedSystem_port_1_cast <= Delay1No185_out;
   Product111_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product111_impl_out,
                 X => Delay1No184_out_to_Product111_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No185_out_to_Product111_impl_parent_implementedSystem_port_1_cast);

SharedReg274_out_to_MUX_Product111_impl_0_parent_implementedSystem_port_1_cast <= SharedReg274_out;
SharedReg309_out_to_MUX_Product111_impl_0_parent_implementedSystem_port_2_cast <= SharedReg309_out;
   MUX_Product111_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg274_out_to_MUX_Product111_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg309_out_to_MUX_Product111_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product111_impl_0_out);

   Delay1No184_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_impl_0_out,
                 Y => Delay1No184_out);

SharedReg75_out_to_MUX_Product111_impl_1_parent_implementedSystem_port_1_cast <= SharedReg75_out;
SharedReg36_out_to_MUX_Product111_impl_1_parent_implementedSystem_port_2_cast <= SharedReg36_out;
   MUX_Product111_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg75_out_to_MUX_Product111_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg36_out_to_MUX_Product111_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product111_impl_1_out);

   Delay1No185_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_impl_1_out,
                 Y => Delay1No185_out);

Delay1No186_out_to_Product210_impl_parent_implementedSystem_port_0_cast <= Delay1No186_out;
Delay1No187_out_to_Product210_impl_parent_implementedSystem_port_1_cast <= Delay1No187_out;
   Product210_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product210_impl_out,
                 X => Delay1No186_out_to_Product210_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No187_out_to_Product210_impl_parent_implementedSystem_port_1_cast);

SharedReg275_out_to_MUX_Product210_impl_0_parent_implementedSystem_port_1_cast <= SharedReg275_out;
SharedReg37_out_to_MUX_Product210_impl_0_parent_implementedSystem_port_2_cast <= SharedReg37_out;
   MUX_Product210_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg275_out_to_MUX_Product210_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg37_out_to_MUX_Product210_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product210_impl_0_out);

   Delay1No186_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_impl_0_out,
                 Y => Delay1No186_out);

SharedReg74_out_to_MUX_Product210_impl_1_parent_implementedSystem_port_1_cast <= SharedReg74_out;
SharedReg309_out_to_MUX_Product210_impl_1_parent_implementedSystem_port_2_cast <= SharedReg309_out;
   MUX_Product210_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg74_out_to_MUX_Product210_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg309_out_to_MUX_Product210_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product210_impl_1_out);

   Delay1No187_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_impl_1_out,
                 Y => Delay1No187_out);

Delay1No188_out_to_Product310_impl_parent_implementedSystem_port_0_cast <= Delay1No188_out;
Delay1No189_out_to_Product310_impl_parent_implementedSystem_port_1_cast <= Delay1No189_out;
   Product310_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product310_impl_out,
                 X => Delay1No188_out_to_Product310_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No189_out_to_Product310_impl_parent_implementedSystem_port_1_cast);

SharedReg75_out_to_MUX_Product310_impl_0_parent_implementedSystem_port_1_cast <= SharedReg75_out;
SharedReg334_out_to_MUX_Product310_impl_0_parent_implementedSystem_port_2_cast <= SharedReg334_out;
   MUX_Product310_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg75_out_to_MUX_Product310_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg334_out_to_MUX_Product310_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product310_impl_0_out);

   Delay1No188_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_impl_0_out,
                 Y => Delay1No188_out);

SharedReg275_out_to_MUX_Product310_impl_1_parent_implementedSystem_port_1_cast <= SharedReg275_out;
SharedReg61_out_to_MUX_Product310_impl_1_parent_implementedSystem_port_2_cast <= SharedReg61_out;
   MUX_Product310_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg275_out_to_MUX_Product310_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg61_out_to_MUX_Product310_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product310_impl_1_out);

   Delay1No189_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_impl_1_out,
                 Y => Delay1No189_out);

Delay1No190_out_to_Subtract11_impl_parent_implementedSystem_port_0_cast <= Delay1No190_out;
Delay1No191_out_to_Subtract11_impl_parent_implementedSystem_port_1_cast <= Delay1No191_out;
   Subtract11_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract11_impl_out,
                 X => Delay1No190_out_to_Subtract11_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No191_out_to_Subtract11_impl_parent_implementedSystem_port_1_cast);

SharedReg119_out_to_MUX_Subtract11_impl_0_parent_implementedSystem_port_1_cast <= SharedReg119_out;
SharedReg97_out_to_MUX_Subtract11_impl_0_parent_implementedSystem_port_2_cast <= SharedReg97_out;
   MUX_Subtract11_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg119_out_to_MUX_Subtract11_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg97_out_to_MUX_Subtract11_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract11_impl_0_out);

   Delay1No190_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract11_impl_0_out,
                 Y => Delay1No190_out);

SharedReg122_out_to_MUX_Subtract11_impl_1_parent_implementedSystem_port_1_cast <= SharedReg122_out;
SharedReg91_out_to_MUX_Subtract11_impl_1_parent_implementedSystem_port_2_cast <= SharedReg91_out;
   MUX_Subtract11_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg122_out_to_MUX_Subtract11_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg91_out_to_MUX_Subtract11_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract11_impl_1_out);

   Delay1No191_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract11_impl_1_out,
                 Y => Delay1No191_out);

Delay1No192_out_to_Add53_impl_parent_implementedSystem_port_0_cast <= Delay1No192_out;
Delay1No193_out_to_Add53_impl_parent_implementedSystem_port_1_cast <= Delay1No193_out;
   Add53_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add53_impl_out,
                 X => Delay1No192_out_to_Add53_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No193_out_to_Add53_impl_parent_implementedSystem_port_1_cast);

SharedReg126_out_to_MUX_Add53_impl_0_parent_implementedSystem_port_1_cast <= SharedReg126_out;
SharedReg98_out_to_MUX_Add53_impl_0_parent_implementedSystem_port_2_cast <= SharedReg98_out;
   MUX_Add53_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg126_out_to_MUX_Add53_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg98_out_to_MUX_Add53_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add53_impl_0_out);

   Delay1No192_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add53_impl_0_out,
                 Y => Delay1No192_out);

SharedReg127_out_to_MUX_Add53_impl_1_parent_implementedSystem_port_1_cast <= SharedReg127_out;
SharedReg88_out_to_MUX_Add53_impl_1_parent_implementedSystem_port_2_cast <= SharedReg88_out;
   MUX_Add53_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg127_out_to_MUX_Add53_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg88_out_to_MUX_Add53_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add53_impl_1_out);

   Delay1No193_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add53_impl_1_out,
                 Y => Delay1No193_out);

Delay1No194_out_to_Product40_impl_parent_implementedSystem_port_0_cast <= Delay1No194_out;
Delay1No195_out_to_Product40_impl_parent_implementedSystem_port_1_cast <= Delay1No195_out;
   Product40_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product40_impl_out,
                 X => Delay1No194_out_to_Product40_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No195_out_to_Product40_impl_parent_implementedSystem_port_1_cast);

SharedReg276_out_to_MUX_Product40_impl_0_parent_implementedSystem_port_1_cast <= SharedReg276_out;
SharedReg334_out_to_MUX_Product40_impl_0_parent_implementedSystem_port_2_cast <= SharedReg334_out;
   MUX_Product40_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg276_out_to_MUX_Product40_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg334_out_to_MUX_Product40_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product40_impl_0_out);

   Delay1No194_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product40_impl_0_out,
                 Y => Delay1No194_out);

SharedReg37_out_to_MUX_Product40_impl_1_parent_implementedSystem_port_1_cast <= SharedReg37_out;
SharedReg63_out_to_MUX_Product40_impl_1_parent_implementedSystem_port_2_cast <= SharedReg63_out;
   MUX_Product40_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg37_out_to_MUX_Product40_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg63_out_to_MUX_Product40_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product40_impl_1_out);

   Delay1No195_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product40_impl_1_out,
                 Y => Delay1No195_out);

Delay1No196_out_to_Product112_impl_parent_implementedSystem_port_0_cast <= Delay1No196_out;
Delay1No197_out_to_Product112_impl_parent_implementedSystem_port_1_cast <= Delay1No197_out;
   Product112_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product112_impl_out,
                 X => Delay1No196_out_to_Product112_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No197_out_to_Product112_impl_parent_implementedSystem_port_1_cast);

SharedReg276_out_to_MUX_Product112_impl_0_parent_implementedSystem_port_1_cast <= SharedReg276_out;
SharedReg335_out_to_MUX_Product112_impl_0_parent_implementedSystem_port_2_cast <= SharedReg335_out;
   MUX_Product112_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg276_out_to_MUX_Product112_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg335_out_to_MUX_Product112_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product112_impl_0_out);

   Delay1No196_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product112_impl_0_out,
                 Y => Delay1No196_out);

SharedReg38_out_to_MUX_Product112_impl_1_parent_implementedSystem_port_1_cast <= SharedReg38_out;
SharedReg61_out_to_MUX_Product112_impl_1_parent_implementedSystem_port_2_cast <= SharedReg61_out;
   MUX_Product112_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg38_out_to_MUX_Product112_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg61_out_to_MUX_Product112_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product112_impl_1_out);

   Delay1No197_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product112_impl_1_out,
                 Y => Delay1No197_out);

Delay1No198_out_to_Product211_impl_parent_implementedSystem_port_0_cast <= Delay1No198_out;
Delay1No199_out_to_Product211_impl_parent_implementedSystem_port_1_cast <= Delay1No199_out;
   Product211_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product211_impl_out,
                 X => Delay1No198_out_to_Product211_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No199_out_to_Product211_impl_parent_implementedSystem_port_1_cast);

SharedReg277_out_to_MUX_Product211_impl_0_parent_implementedSystem_port_1_cast <= SharedReg277_out;
SharedReg63_out_to_MUX_Product211_impl_0_parent_implementedSystem_port_2_cast <= SharedReg63_out;
   MUX_Product211_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg277_out_to_MUX_Product211_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg63_out_to_MUX_Product211_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product211_impl_0_out);

   Delay1No198_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product211_impl_0_out,
                 Y => Delay1No198_out);

SharedReg37_out_to_MUX_Product211_impl_1_parent_implementedSystem_port_1_cast <= SharedReg37_out;
SharedReg335_out_to_MUX_Product211_impl_1_parent_implementedSystem_port_2_cast <= SharedReg335_out;
   MUX_Product211_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg37_out_to_MUX_Product211_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg335_out_to_MUX_Product211_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product211_impl_1_out);

   Delay1No199_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product211_impl_1_out,
                 Y => Delay1No199_out);

Delay1No200_out_to_Product311_impl_parent_implementedSystem_port_0_cast <= Delay1No200_out;
Delay1No201_out_to_Product311_impl_parent_implementedSystem_port_1_cast <= Delay1No201_out;
   Product311_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product311_impl_out,
                 X => Delay1No200_out_to_Product311_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No201_out_to_Product311_impl_parent_implementedSystem_port_1_cast);

SharedReg38_out_to_MUX_Product311_impl_0_parent_implementedSystem_port_1_cast <= SharedReg38_out;
SharedReg47_out_to_MUX_Product311_impl_0_parent_implementedSystem_port_2_cast <= SharedReg47_out;
   MUX_Product311_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg38_out_to_MUX_Product311_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg47_out_to_MUX_Product311_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product311_impl_0_out);

   Delay1No200_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product311_impl_0_out,
                 Y => Delay1No200_out);

SharedReg277_out_to_MUX_Product311_impl_1_parent_implementedSystem_port_1_cast <= SharedReg277_out;
SharedReg311_out_to_MUX_Product311_impl_1_parent_implementedSystem_port_2_cast <= SharedReg311_out;
   MUX_Product311_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg277_out_to_MUX_Product311_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg311_out_to_MUX_Product311_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product311_impl_1_out);

   Delay1No201_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product311_impl_1_out,
                 Y => Delay1No201_out);

Delay1No202_out_to_Subtract12_impl_parent_implementedSystem_port_0_cast <= Delay1No202_out;
Delay1No203_out_to_Subtract12_impl_parent_implementedSystem_port_1_cast <= Delay1No203_out;
   Subtract12_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract12_impl_out,
                 X => Delay1No202_out_to_Subtract12_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No203_out_to_Subtract12_impl_parent_implementedSystem_port_1_cast);

SharedReg125_out_to_MUX_Subtract12_impl_0_parent_implementedSystem_port_1_cast <= SharedReg125_out;
SharedReg131_out_to_MUX_Subtract12_impl_0_parent_implementedSystem_port_2_cast <= SharedReg131_out;
   MUX_Subtract12_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg125_out_to_MUX_Subtract12_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg131_out_to_MUX_Subtract12_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract12_impl_0_out);

   Delay1No202_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_impl_0_out,
                 Y => Delay1No202_out);

SharedReg128_out_to_MUX_Subtract12_impl_1_parent_implementedSystem_port_1_cast <= SharedReg128_out;
SharedReg134_out_to_MUX_Subtract12_impl_1_parent_implementedSystem_port_2_cast <= SharedReg134_out;
   MUX_Subtract12_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg128_out_to_MUX_Subtract12_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg134_out_to_MUX_Subtract12_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract12_impl_1_out);

   Delay1No203_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_impl_1_out,
                 Y => Delay1No203_out);

Delay1No204_out_to_Add54_impl_parent_implementedSystem_port_0_cast <= Delay1No204_out;
Delay1No205_out_to_Add54_impl_parent_implementedSystem_port_1_cast <= Delay1No205_out;
   Add54_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add54_impl_out,
                 X => Delay1No204_out_to_Add54_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No205_out_to_Add54_impl_parent_implementedSystem_port_1_cast);

SharedReg132_out_to_MUX_Add54_impl_0_parent_implementedSystem_port_1_cast <= SharedReg132_out;
SharedReg138_out_to_MUX_Add54_impl_0_parent_implementedSystem_port_2_cast <= SharedReg138_out;
   MUX_Add54_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg132_out_to_MUX_Add54_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg138_out_to_MUX_Add54_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add54_impl_0_out);

   Delay1No204_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add54_impl_0_out,
                 Y => Delay1No204_out);

SharedReg133_out_to_MUX_Add54_impl_1_parent_implementedSystem_port_1_cast <= SharedReg133_out;
SharedReg139_out_to_MUX_Add54_impl_1_parent_implementedSystem_port_2_cast <= SharedReg139_out;
   MUX_Add54_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg133_out_to_MUX_Add54_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg139_out_to_MUX_Add54_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add54_impl_1_out);

   Delay1No205_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add54_impl_1_out,
                 Y => Delay1No205_out);

Delay1No206_out_to_Product41_impl_parent_implementedSystem_port_0_cast <= Delay1No206_out;
Delay1No207_out_to_Product41_impl_parent_implementedSystem_port_1_cast <= Delay1No207_out;
   Product41_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product41_impl_out,
                 X => Delay1No206_out_to_Product41_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No207_out_to_Product41_impl_parent_implementedSystem_port_1_cast);

SharedReg278_out_to_MUX_Product41_impl_0_parent_implementedSystem_port_1_cast <= SharedReg278_out;
SharedReg314_out_to_MUX_Product41_impl_0_parent_implementedSystem_port_2_cast <= SharedReg314_out;
   MUX_Product41_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg278_out_to_MUX_Product41_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg314_out_to_MUX_Product41_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product41_impl_0_out);

   Delay1No206_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product41_impl_0_out,
                 Y => Delay1No206_out);

SharedReg39_out_to_MUX_Product41_impl_1_parent_implementedSystem_port_1_cast <= SharedReg39_out;
SharedReg38_out_to_MUX_Product41_impl_1_parent_implementedSystem_port_2_cast <= SharedReg38_out;
   MUX_Product41_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg39_out_to_MUX_Product41_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg38_out_to_MUX_Product41_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product41_impl_1_out);

   Delay1No207_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product41_impl_1_out,
                 Y => Delay1No207_out);

Delay1No208_out_to_Product113_impl_parent_implementedSystem_port_0_cast <= Delay1No208_out;
Delay1No209_out_to_Product113_impl_parent_implementedSystem_port_1_cast <= Delay1No209_out;
   Product113_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product113_impl_out,
                 X => Delay1No208_out_to_Product113_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No209_out_to_Product113_impl_parent_implementedSystem_port_1_cast);

SharedReg278_out_to_MUX_Product113_impl_0_parent_implementedSystem_port_1_cast <= SharedReg278_out;
SharedReg314_out_to_MUX_Product113_impl_0_parent_implementedSystem_port_2_cast <= SharedReg314_out;
   MUX_Product113_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg278_out_to_MUX_Product113_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg314_out_to_MUX_Product113_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product113_impl_0_out);

   Delay1No208_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product113_impl_0_out,
                 Y => Delay1No208_out);

SharedReg40_out_to_MUX_Product113_impl_1_parent_implementedSystem_port_1_cast <= SharedReg40_out;
SharedReg39_out_to_MUX_Product113_impl_1_parent_implementedSystem_port_2_cast <= SharedReg39_out;
   MUX_Product113_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg40_out_to_MUX_Product113_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg39_out_to_MUX_Product113_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product113_impl_1_out);

   Delay1No209_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product113_impl_1_out,
                 Y => Delay1No209_out);

Delay1No210_out_to_Product212_impl_parent_implementedSystem_port_0_cast <= Delay1No210_out;
Delay1No211_out_to_Product212_impl_parent_implementedSystem_port_1_cast <= Delay1No211_out;
   Product212_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product212_impl_out,
                 X => Delay1No210_out_to_Product212_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No211_out_to_Product212_impl_parent_implementedSystem_port_1_cast);

SharedReg279_out_to_MUX_Product212_impl_0_parent_implementedSystem_port_1_cast <= SharedReg279_out;
SharedReg315_out_to_MUX_Product212_impl_0_parent_implementedSystem_port_2_cast <= SharedReg315_out;
   MUX_Product212_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg279_out_to_MUX_Product212_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg315_out_to_MUX_Product212_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product212_impl_0_out);

   Delay1No210_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product212_impl_0_out,
                 Y => Delay1No210_out);

SharedReg39_out_to_MUX_Product212_impl_1_parent_implementedSystem_port_1_cast <= SharedReg39_out;
SharedReg38_out_to_MUX_Product212_impl_1_parent_implementedSystem_port_2_cast <= SharedReg38_out;
   MUX_Product212_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg39_out_to_MUX_Product212_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg38_out_to_MUX_Product212_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product212_impl_1_out);

   Delay1No211_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product212_impl_1_out,
                 Y => Delay1No211_out);

Delay1No212_out_to_Product312_impl_parent_implementedSystem_port_0_cast <= Delay1No212_out;
Delay1No213_out_to_Product312_impl_parent_implementedSystem_port_1_cast <= Delay1No213_out;
   Product312_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product312_impl_out,
                 X => Delay1No212_out_to_Product312_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No213_out_to_Product312_impl_parent_implementedSystem_port_1_cast);

SharedReg40_out_to_MUX_Product312_impl_0_parent_implementedSystem_port_1_cast <= SharedReg40_out;
SharedReg39_out_to_MUX_Product312_impl_0_parent_implementedSystem_port_2_cast <= SharedReg39_out;
   MUX_Product312_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg40_out_to_MUX_Product312_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg39_out_to_MUX_Product312_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product312_impl_0_out);

   Delay1No212_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product312_impl_0_out,
                 Y => Delay1No212_out);

SharedReg279_out_to_MUX_Product312_impl_1_parent_implementedSystem_port_1_cast <= SharedReg279_out;
SharedReg315_out_to_MUX_Product312_impl_1_parent_implementedSystem_port_2_cast <= SharedReg315_out;
   MUX_Product312_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg279_out_to_MUX_Product312_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg315_out_to_MUX_Product312_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product312_impl_1_out);

   Delay1No213_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product312_impl_1_out,
                 Y => Delay1No213_out);

Delay1No214_out_to_Subtract13_impl_parent_implementedSystem_port_0_cast <= Delay1No214_out;
Delay1No215_out_to_Subtract13_impl_parent_implementedSystem_port_1_cast <= Delay1No215_out;
   Subtract13_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract13_impl_out,
                 X => Delay1No214_out_to_Subtract13_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No215_out_to_Subtract13_impl_parent_implementedSystem_port_1_cast);

SharedReg131_out_to_MUX_Subtract13_impl_0_parent_implementedSystem_port_1_cast <= SharedReg131_out;
SharedReg137_out_to_MUX_Subtract13_impl_0_parent_implementedSystem_port_2_cast <= SharedReg137_out;
   MUX_Subtract13_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg131_out_to_MUX_Subtract13_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg137_out_to_MUX_Subtract13_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract13_impl_0_out);

   Delay1No214_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract13_impl_0_out,
                 Y => Delay1No214_out);

SharedReg134_out_to_MUX_Subtract13_impl_1_parent_implementedSystem_port_1_cast <= SharedReg134_out;
SharedReg140_out_to_MUX_Subtract13_impl_1_parent_implementedSystem_port_2_cast <= SharedReg140_out;
   MUX_Subtract13_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg134_out_to_MUX_Subtract13_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg140_out_to_MUX_Subtract13_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract13_impl_1_out);

   Delay1No215_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract13_impl_1_out,
                 Y => Delay1No215_out);

Delay1No216_out_to_Add56_impl_parent_implementedSystem_port_0_cast <= Delay1No216_out;
Delay1No217_out_to_Add56_impl_parent_implementedSystem_port_1_cast <= Delay1No217_out;
   Add56_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add56_impl_out,
                 X => Delay1No216_out_to_Add56_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No217_out_to_Add56_impl_parent_implementedSystem_port_1_cast);

SharedReg138_out_to_MUX_Add56_impl_0_parent_implementedSystem_port_1_cast <= SharedReg138_out;
SharedReg144_out_to_MUX_Add56_impl_0_parent_implementedSystem_port_2_cast <= SharedReg144_out;
   MUX_Add56_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg138_out_to_MUX_Add56_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg144_out_to_MUX_Add56_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add56_impl_0_out);

   Delay1No216_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add56_impl_0_out,
                 Y => Delay1No216_out);

SharedReg139_out_to_MUX_Add56_impl_1_parent_implementedSystem_port_1_cast <= SharedReg139_out;
SharedReg145_out_to_MUX_Add56_impl_1_parent_implementedSystem_port_2_cast <= SharedReg145_out;
   MUX_Add56_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg139_out_to_MUX_Add56_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg145_out_to_MUX_Add56_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add56_impl_1_out);

   Delay1No217_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add56_impl_1_out,
                 Y => Delay1No217_out);

Delay1No218_out_to_Product43_impl_parent_implementedSystem_port_0_cast <= Delay1No218_out;
Delay1No219_out_to_Product43_impl_parent_implementedSystem_port_1_cast <= Delay1No219_out;
   Product43_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product43_impl_out,
                 X => Delay1No218_out_to_Product43_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No219_out_to_Product43_impl_parent_implementedSystem_port_1_cast);

SharedReg282_out_to_MUX_Product43_impl_0_parent_implementedSystem_port_1_cast <= SharedReg282_out;
SharedReg316_out_to_MUX_Product43_impl_0_parent_implementedSystem_port_2_cast <= SharedReg316_out;
   MUX_Product43_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg282_out_to_MUX_Product43_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg316_out_to_MUX_Product43_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product43_impl_0_out);

   Delay1No218_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product43_impl_0_out,
                 Y => Delay1No218_out);

SharedReg41_out_to_MUX_Product43_impl_1_parent_implementedSystem_port_1_cast <= SharedReg41_out;
SharedReg49_out_to_MUX_Product43_impl_1_parent_implementedSystem_port_2_cast <= SharedReg49_out;
   MUX_Product43_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg41_out_to_MUX_Product43_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg49_out_to_MUX_Product43_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product43_impl_1_out);

   Delay1No219_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product43_impl_1_out,
                 Y => Delay1No219_out);

Delay1No220_out_to_Product115_impl_parent_implementedSystem_port_0_cast <= Delay1No220_out;
Delay1No221_out_to_Product115_impl_parent_implementedSystem_port_1_cast <= Delay1No221_out;
   Product115_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product115_impl_out,
                 X => Delay1No220_out_to_Product115_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No221_out_to_Product115_impl_parent_implementedSystem_port_1_cast);

SharedReg282_out_to_MUX_Product115_impl_0_parent_implementedSystem_port_1_cast <= SharedReg282_out;
SharedReg316_out_to_MUX_Product115_impl_0_parent_implementedSystem_port_2_cast <= SharedReg316_out;
   MUX_Product115_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg282_out_to_MUX_Product115_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg316_out_to_MUX_Product115_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product115_impl_0_out);

   Delay1No220_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product115_impl_0_out,
                 Y => Delay1No220_out);

SharedReg32_out_to_MUX_Product115_impl_1_parent_implementedSystem_port_1_cast <= SharedReg32_out;
SharedReg51_out_to_MUX_Product115_impl_1_parent_implementedSystem_port_2_cast <= SharedReg51_out;
   MUX_Product115_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg32_out_to_MUX_Product115_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg51_out_to_MUX_Product115_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product115_impl_1_out);

   Delay1No221_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product115_impl_1_out,
                 Y => Delay1No221_out);

Delay1No222_out_to_Product214_impl_parent_implementedSystem_port_0_cast <= Delay1No222_out;
Delay1No223_out_to_Product214_impl_parent_implementedSystem_port_1_cast <= Delay1No223_out;
   Product214_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product214_impl_out,
                 X => Delay1No222_out_to_Product214_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No223_out_to_Product214_impl_parent_implementedSystem_port_1_cast);

SharedReg283_out_to_MUX_Product214_impl_0_parent_implementedSystem_port_1_cast <= SharedReg283_out;
SharedReg317_out_to_MUX_Product214_impl_0_parent_implementedSystem_port_2_cast <= SharedReg317_out;
   MUX_Product214_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg283_out_to_MUX_Product214_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg317_out_to_MUX_Product214_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product214_impl_0_out);

   Delay1No222_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product214_impl_0_out,
                 Y => Delay1No222_out);

SharedReg41_out_to_MUX_Product214_impl_1_parent_implementedSystem_port_1_cast <= SharedReg41_out;
SharedReg49_out_to_MUX_Product214_impl_1_parent_implementedSystem_port_2_cast <= SharedReg49_out;
   MUX_Product214_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg41_out_to_MUX_Product214_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg49_out_to_MUX_Product214_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product214_impl_1_out);

   Delay1No223_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product214_impl_1_out,
                 Y => Delay1No223_out);

Delay1No224_out_to_Product314_impl_parent_implementedSystem_port_0_cast <= Delay1No224_out;
Delay1No225_out_to_Product314_impl_parent_implementedSystem_port_1_cast <= Delay1No225_out;
   Product314_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product314_impl_out,
                 X => Delay1No224_out_to_Product314_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No225_out_to_Product314_impl_parent_implementedSystem_port_1_cast);

SharedReg32_out_to_MUX_Product314_impl_0_parent_implementedSystem_port_1_cast <= SharedReg32_out;
SharedReg51_out_to_MUX_Product314_impl_0_parent_implementedSystem_port_2_cast <= SharedReg51_out;
   MUX_Product314_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg32_out_to_MUX_Product314_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg51_out_to_MUX_Product314_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product314_impl_0_out);

   Delay1No224_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product314_impl_0_out,
                 Y => Delay1No224_out);

SharedReg283_out_to_MUX_Product314_impl_1_parent_implementedSystem_port_1_cast <= SharedReg283_out;
SharedReg317_out_to_MUX_Product314_impl_1_parent_implementedSystem_port_2_cast <= SharedReg317_out;
   MUX_Product314_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg283_out_to_MUX_Product314_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg317_out_to_MUX_Product314_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product314_impl_1_out);

   Delay1No225_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product314_impl_1_out,
                 Y => Delay1No225_out);

Delay1No226_out_to_Subtract15_impl_parent_implementedSystem_port_0_cast <= Delay1No226_out;
Delay1No227_out_to_Subtract15_impl_parent_implementedSystem_port_1_cast <= Delay1No227_out;
   Subtract15_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract15_impl_out,
                 X => Delay1No226_out_to_Subtract15_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No227_out_to_Subtract15_impl_parent_implementedSystem_port_1_cast);

SharedReg137_out_to_MUX_Subtract15_impl_0_parent_implementedSystem_port_1_cast <= SharedReg137_out;
SharedReg143_out_to_MUX_Subtract15_impl_0_parent_implementedSystem_port_2_cast <= SharedReg143_out;
   MUX_Subtract15_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg137_out_to_MUX_Subtract15_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg143_out_to_MUX_Subtract15_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract15_impl_0_out);

   Delay1No226_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract15_impl_0_out,
                 Y => Delay1No226_out);

SharedReg140_out_to_MUX_Subtract15_impl_1_parent_implementedSystem_port_1_cast <= SharedReg140_out;
SharedReg146_out_to_MUX_Subtract15_impl_1_parent_implementedSystem_port_2_cast <= SharedReg146_out;
   MUX_Subtract15_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg140_out_to_MUX_Subtract15_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg146_out_to_MUX_Subtract15_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract15_impl_1_out);

   Delay1No227_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract15_impl_1_out,
                 Y => Delay1No227_out);

Delay1No228_out_to_Add57_impl_parent_implementedSystem_port_0_cast <= Delay1No228_out;
Delay1No229_out_to_Add57_impl_parent_implementedSystem_port_1_cast <= Delay1No229_out;
   Add57_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add57_impl_out,
                 X => Delay1No228_out_to_Add57_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No229_out_to_Add57_impl_parent_implementedSystem_port_1_cast);

SharedReg144_out_to_MUX_Add57_impl_0_parent_implementedSystem_port_1_cast <= SharedReg144_out;
SharedReg150_out_to_MUX_Add57_impl_0_parent_implementedSystem_port_2_cast <= SharedReg150_out;
   MUX_Add57_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg144_out_to_MUX_Add57_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg150_out_to_MUX_Add57_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add57_impl_0_out);

   Delay1No228_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add57_impl_0_out,
                 Y => Delay1No228_out);

SharedReg145_out_to_MUX_Add57_impl_1_parent_implementedSystem_port_1_cast <= SharedReg145_out;
SharedReg151_out_to_MUX_Add57_impl_1_parent_implementedSystem_port_2_cast <= SharedReg151_out;
   MUX_Add57_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg145_out_to_MUX_Add57_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg151_out_to_MUX_Add57_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add57_impl_1_out);

   Delay1No229_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add57_impl_1_out,
                 Y => Delay1No229_out);

Delay1No230_out_to_Product44_impl_parent_implementedSystem_port_0_cast <= Delay1No230_out;
Delay1No231_out_to_Product44_impl_parent_implementedSystem_port_1_cast <= Delay1No231_out;
   Product44_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product44_impl_out,
                 X => Delay1No230_out_to_Product44_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No231_out_to_Product44_impl_parent_implementedSystem_port_1_cast);

SharedReg284_out_to_MUX_Product44_impl_0_parent_implementedSystem_port_1_cast <= SharedReg284_out;
SharedReg320_out_to_MUX_Product44_impl_0_parent_implementedSystem_port_2_cast <= SharedReg320_out;
   MUX_Product44_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg284_out_to_MUX_Product44_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg320_out_to_MUX_Product44_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product44_impl_0_out);

   Delay1No230_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product44_impl_0_out,
                 Y => Delay1No230_out);

SharedReg42_out_to_MUX_Product44_impl_1_parent_implementedSystem_port_1_cast <= SharedReg42_out;
SharedReg229_out_to_MUX_Product44_impl_1_parent_implementedSystem_port_2_cast <= SharedReg229_out;
   MUX_Product44_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg42_out_to_MUX_Product44_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg229_out_to_MUX_Product44_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product44_impl_1_out);

   Delay1No231_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product44_impl_1_out,
                 Y => Delay1No231_out);

Delay1No232_out_to_Product116_impl_parent_implementedSystem_port_0_cast <= Delay1No232_out;
Delay1No233_out_to_Product116_impl_parent_implementedSystem_port_1_cast <= Delay1No233_out;
   Product116_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product116_impl_out,
                 X => Delay1No232_out_to_Product116_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No233_out_to_Product116_impl_parent_implementedSystem_port_1_cast);

SharedReg284_out_to_MUX_Product116_impl_0_parent_implementedSystem_port_1_cast <= SharedReg284_out;
SharedReg320_out_to_MUX_Product116_impl_0_parent_implementedSystem_port_2_cast <= SharedReg320_out;
   MUX_Product116_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg284_out_to_MUX_Product116_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg320_out_to_MUX_Product116_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product116_impl_0_out);

   Delay1No232_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product116_impl_0_out,
                 Y => Delay1No232_out);

SharedReg43_out_to_MUX_Product116_impl_1_parent_implementedSystem_port_1_cast <= SharedReg43_out;
SharedReg230_out_to_MUX_Product116_impl_1_parent_implementedSystem_port_2_cast <= SharedReg230_out;
   MUX_Product116_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg43_out_to_MUX_Product116_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg230_out_to_MUX_Product116_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product116_impl_1_out);

   Delay1No233_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product116_impl_1_out,
                 Y => Delay1No233_out);

Delay1No234_out_to_Product215_impl_parent_implementedSystem_port_0_cast <= Delay1No234_out;
Delay1No235_out_to_Product215_impl_parent_implementedSystem_port_1_cast <= Delay1No235_out;
   Product215_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product215_impl_out,
                 X => Delay1No234_out_to_Product215_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No235_out_to_Product215_impl_parent_implementedSystem_port_1_cast);

SharedReg285_out_to_MUX_Product215_impl_0_parent_implementedSystem_port_1_cast <= SharedReg285_out;
SharedReg321_out_to_MUX_Product215_impl_0_parent_implementedSystem_port_2_cast <= SharedReg321_out;
   MUX_Product215_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg285_out_to_MUX_Product215_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg321_out_to_MUX_Product215_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product215_impl_0_out);

   Delay1No234_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product215_impl_0_out,
                 Y => Delay1No234_out);

SharedReg42_out_to_MUX_Product215_impl_1_parent_implementedSystem_port_1_cast <= SharedReg42_out;
SharedReg229_out_to_MUX_Product215_impl_1_parent_implementedSystem_port_2_cast <= SharedReg229_out;
   MUX_Product215_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg42_out_to_MUX_Product215_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg229_out_to_MUX_Product215_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product215_impl_1_out);

   Delay1No235_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product215_impl_1_out,
                 Y => Delay1No235_out);

Delay1No236_out_to_Product315_impl_parent_implementedSystem_port_0_cast <= Delay1No236_out;
Delay1No237_out_to_Product315_impl_parent_implementedSystem_port_1_cast <= Delay1No237_out;
   Product315_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product315_impl_out,
                 X => Delay1No236_out_to_Product315_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No237_out_to_Product315_impl_parent_implementedSystem_port_1_cast);

SharedReg43_out_to_MUX_Product315_impl_0_parent_implementedSystem_port_1_cast <= SharedReg43_out;
SharedReg230_out_to_MUX_Product315_impl_0_parent_implementedSystem_port_2_cast <= SharedReg230_out;
   MUX_Product315_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg43_out_to_MUX_Product315_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg230_out_to_MUX_Product315_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product315_impl_0_out);

   Delay1No236_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product315_impl_0_out,
                 Y => Delay1No236_out);

SharedReg285_out_to_MUX_Product315_impl_1_parent_implementedSystem_port_1_cast <= SharedReg285_out;
SharedReg321_out_to_MUX_Product315_impl_1_parent_implementedSystem_port_2_cast <= SharedReg321_out;
   MUX_Product315_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg285_out_to_MUX_Product315_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg321_out_to_MUX_Product315_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product315_impl_1_out);

   Delay1No237_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product315_impl_1_out,
                 Y => Delay1No237_out);

Delay1No238_out_to_Subtract16_impl_parent_implementedSystem_port_0_cast <= Delay1No238_out;
Delay1No239_out_to_Subtract16_impl_parent_implementedSystem_port_1_cast <= Delay1No239_out;
   Subtract16_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract16_impl_out,
                 X => Delay1No238_out_to_Subtract16_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No239_out_to_Subtract16_impl_parent_implementedSystem_port_1_cast);

SharedReg143_out_to_MUX_Subtract16_impl_0_parent_implementedSystem_port_1_cast <= SharedReg143_out;
SharedReg149_out_to_MUX_Subtract16_impl_0_parent_implementedSystem_port_2_cast <= SharedReg149_out;
   MUX_Subtract16_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg143_out_to_MUX_Subtract16_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg149_out_to_MUX_Subtract16_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract16_impl_0_out);

   Delay1No238_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract16_impl_0_out,
                 Y => Delay1No238_out);

SharedReg146_out_to_MUX_Subtract16_impl_1_parent_implementedSystem_port_1_cast <= SharedReg146_out;
SharedReg152_out_to_MUX_Subtract16_impl_1_parent_implementedSystem_port_2_cast <= SharedReg152_out;
   MUX_Subtract16_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg146_out_to_MUX_Subtract16_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg152_out_to_MUX_Subtract16_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract16_impl_1_out);

   Delay1No239_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract16_impl_1_out,
                 Y => Delay1No239_out);

Delay1No240_out_to_Add58_impl_parent_implementedSystem_port_0_cast <= Delay1No240_out;
Delay1No241_out_to_Add58_impl_parent_implementedSystem_port_1_cast <= Delay1No241_out;
   Add58_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add58_impl_out,
                 X => Delay1No240_out_to_Add58_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No241_out_to_Add58_impl_parent_implementedSystem_port_1_cast);

SharedReg150_out_to_MUX_Add58_impl_0_parent_implementedSystem_port_1_cast <= SharedReg150_out;
SharedReg156_out_to_MUX_Add58_impl_0_parent_implementedSystem_port_2_cast <= SharedReg156_out;
   MUX_Add58_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg150_out_to_MUX_Add58_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg156_out_to_MUX_Add58_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add58_impl_0_out);

   Delay1No240_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add58_impl_0_out,
                 Y => Delay1No240_out);

SharedReg151_out_to_MUX_Add58_impl_1_parent_implementedSystem_port_1_cast <= SharedReg151_out;
SharedReg157_out_to_MUX_Add58_impl_1_parent_implementedSystem_port_2_cast <= SharedReg157_out;
   MUX_Add58_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg151_out_to_MUX_Add58_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg157_out_to_MUX_Add58_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add58_impl_1_out);

   Delay1No241_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add58_impl_1_out,
                 Y => Delay1No241_out);

Delay1No242_out_to_Product45_impl_parent_implementedSystem_port_0_cast <= Delay1No242_out;
Delay1No243_out_to_Product45_impl_parent_implementedSystem_port_1_cast <= Delay1No243_out;
   Product45_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product45_impl_out,
                 X => Delay1No242_out_to_Product45_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No243_out_to_Product45_impl_parent_implementedSystem_port_1_cast);

SharedReg286_out_to_MUX_Product45_impl_0_parent_implementedSystem_port_1_cast <= SharedReg286_out;
SharedReg318_out_to_MUX_Product45_impl_0_parent_implementedSystem_port_2_cast <= SharedReg318_out;
   MUX_Product45_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg286_out_to_MUX_Product45_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg318_out_to_MUX_Product45_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product45_impl_0_out);

   Delay1No242_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product45_impl_0_out,
                 Y => Delay1No242_out);

SharedReg226_out_to_MUX_Product45_impl_1_parent_implementedSystem_port_1_cast <= SharedReg226_out;
SharedReg231_out_to_MUX_Product45_impl_1_parent_implementedSystem_port_2_cast <= SharedReg231_out;
   MUX_Product45_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg226_out_to_MUX_Product45_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg231_out_to_MUX_Product45_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product45_impl_1_out);

   Delay1No243_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product45_impl_1_out,
                 Y => Delay1No243_out);

Delay1No244_out_to_Product117_impl_parent_implementedSystem_port_0_cast <= Delay1No244_out;
Delay1No245_out_to_Product117_impl_parent_implementedSystem_port_1_cast <= Delay1No245_out;
   Product117_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product117_impl_out,
                 X => Delay1No244_out_to_Product117_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No245_out_to_Product117_impl_parent_implementedSystem_port_1_cast);

SharedReg286_out_to_MUX_Product117_impl_0_parent_implementedSystem_port_1_cast <= SharedReg286_out;
SharedReg318_out_to_MUX_Product117_impl_0_parent_implementedSystem_port_2_cast <= SharedReg318_out;
   MUX_Product117_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg286_out_to_MUX_Product117_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg318_out_to_MUX_Product117_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product117_impl_0_out);

   Delay1No244_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product117_impl_0_out,
                 Y => Delay1No244_out);

SharedReg227_out_to_MUX_Product117_impl_1_parent_implementedSystem_port_1_cast <= SharedReg227_out;
SharedReg232_out_to_MUX_Product117_impl_1_parent_implementedSystem_port_2_cast <= SharedReg232_out;
   MUX_Product117_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg227_out_to_MUX_Product117_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg232_out_to_MUX_Product117_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product117_impl_1_out);

   Delay1No245_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product117_impl_1_out,
                 Y => Delay1No245_out);

Delay1No246_out_to_Product216_impl_parent_implementedSystem_port_0_cast <= Delay1No246_out;
Delay1No247_out_to_Product216_impl_parent_implementedSystem_port_1_cast <= Delay1No247_out;
   Product216_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product216_impl_out,
                 X => Delay1No246_out_to_Product216_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No247_out_to_Product216_impl_parent_implementedSystem_port_1_cast);

SharedReg287_out_to_MUX_Product216_impl_0_parent_implementedSystem_port_1_cast <= SharedReg287_out;
SharedReg319_out_to_MUX_Product216_impl_0_parent_implementedSystem_port_2_cast <= SharedReg319_out;
   MUX_Product216_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg287_out_to_MUX_Product216_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg319_out_to_MUX_Product216_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product216_impl_0_out);

   Delay1No246_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product216_impl_0_out,
                 Y => Delay1No246_out);

SharedReg226_out_to_MUX_Product216_impl_1_parent_implementedSystem_port_1_cast <= SharedReg226_out;
SharedReg231_out_to_MUX_Product216_impl_1_parent_implementedSystem_port_2_cast <= SharedReg231_out;
   MUX_Product216_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg226_out_to_MUX_Product216_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg231_out_to_MUX_Product216_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product216_impl_1_out);

   Delay1No247_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product216_impl_1_out,
                 Y => Delay1No247_out);

Delay1No248_out_to_Product316_impl_parent_implementedSystem_port_0_cast <= Delay1No248_out;
Delay1No249_out_to_Product316_impl_parent_implementedSystem_port_1_cast <= Delay1No249_out;
   Product316_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product316_impl_out,
                 X => Delay1No248_out_to_Product316_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No249_out_to_Product316_impl_parent_implementedSystem_port_1_cast);

SharedReg227_out_to_MUX_Product316_impl_0_parent_implementedSystem_port_1_cast <= SharedReg227_out;
SharedReg232_out_to_MUX_Product316_impl_0_parent_implementedSystem_port_2_cast <= SharedReg232_out;
   MUX_Product316_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg227_out_to_MUX_Product316_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg232_out_to_MUX_Product316_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product316_impl_0_out);

   Delay1No248_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product316_impl_0_out,
                 Y => Delay1No248_out);

SharedReg287_out_to_MUX_Product316_impl_1_parent_implementedSystem_port_1_cast <= SharedReg287_out;
SharedReg319_out_to_MUX_Product316_impl_1_parent_implementedSystem_port_2_cast <= SharedReg319_out;
   MUX_Product316_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg287_out_to_MUX_Product316_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg319_out_to_MUX_Product316_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product316_impl_1_out);

   Delay1No249_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product316_impl_1_out,
                 Y => Delay1No249_out);

Delay1No250_out_to_Subtract17_impl_parent_implementedSystem_port_0_cast <= Delay1No250_out;
Delay1No251_out_to_Subtract17_impl_parent_implementedSystem_port_1_cast <= Delay1No251_out;
   Subtract17_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract17_impl_out,
                 X => Delay1No250_out_to_Subtract17_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No251_out_to_Subtract17_impl_parent_implementedSystem_port_1_cast);

SharedReg149_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_1_cast <= SharedReg149_out;
SharedReg155_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_2_cast <= SharedReg155_out;
   MUX_Subtract17_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg149_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg155_out_to_MUX_Subtract17_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract17_impl_0_out);

   Delay1No250_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract17_impl_0_out,
                 Y => Delay1No250_out);

SharedReg152_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_1_cast <= SharedReg152_out;
SharedReg158_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_2_cast <= SharedReg158_out;
   MUX_Subtract17_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg152_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg158_out_to_MUX_Subtract17_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract17_impl_1_out);

   Delay1No251_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract17_impl_1_out,
                 Y => Delay1No251_out);

Delay1No252_out_to_Add59_impl_parent_implementedSystem_port_0_cast <= Delay1No252_out;
Delay1No253_out_to_Add59_impl_parent_implementedSystem_port_1_cast <= Delay1No253_out;
   Add59_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add59_impl_out,
                 X => Delay1No252_out_to_Add59_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No253_out_to_Add59_impl_parent_implementedSystem_port_1_cast);

SharedReg156_out_to_MUX_Add59_impl_0_parent_implementedSystem_port_1_cast <= SharedReg156_out;
SharedReg162_out_to_MUX_Add59_impl_0_parent_implementedSystem_port_2_cast <= SharedReg162_out;
   MUX_Add59_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg156_out_to_MUX_Add59_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg162_out_to_MUX_Add59_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add59_impl_0_out);

   Delay1No252_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add59_impl_0_out,
                 Y => Delay1No252_out);

SharedReg157_out_to_MUX_Add59_impl_1_parent_implementedSystem_port_1_cast <= SharedReg157_out;
SharedReg163_out_to_MUX_Add59_impl_1_parent_implementedSystem_port_2_cast <= SharedReg163_out;
   MUX_Add59_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg157_out_to_MUX_Add59_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg163_out_to_MUX_Add59_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add59_impl_1_out);

   Delay1No253_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add59_impl_1_out,
                 Y => Delay1No253_out);

Delay1No254_out_to_Product46_impl_parent_implementedSystem_port_0_cast <= Delay1No254_out;
Delay1No255_out_to_Product46_impl_parent_implementedSystem_port_1_cast <= Delay1No255_out;
   Product46_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product46_impl_out,
                 X => Delay1No254_out_to_Product46_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No255_out_to_Product46_impl_parent_implementedSystem_port_1_cast);

SharedReg288_out_to_MUX_Product46_impl_0_parent_implementedSystem_port_1_cast <= SharedReg288_out;
SharedReg322_out_to_MUX_Product46_impl_0_parent_implementedSystem_port_2_cast <= SharedReg322_out;
   MUX_Product46_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg288_out_to_MUX_Product46_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg322_out_to_MUX_Product46_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product46_impl_0_out);

   Delay1No254_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product46_impl_0_out,
                 Y => Delay1No254_out);

SharedReg228_out_to_MUX_Product46_impl_1_parent_implementedSystem_port_1_cast <= SharedReg228_out;
SharedReg53_out_to_MUX_Product46_impl_1_parent_implementedSystem_port_2_cast <= SharedReg53_out;
   MUX_Product46_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg228_out_to_MUX_Product46_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg53_out_to_MUX_Product46_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product46_impl_1_out);

   Delay1No255_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product46_impl_1_out,
                 Y => Delay1No255_out);

Delay1No256_out_to_Product118_impl_parent_implementedSystem_port_0_cast <= Delay1No256_out;
Delay1No257_out_to_Product118_impl_parent_implementedSystem_port_1_cast <= Delay1No257_out;
   Product118_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product118_impl_out,
                 X => Delay1No256_out_to_Product118_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No257_out_to_Product118_impl_parent_implementedSystem_port_1_cast);

SharedReg288_out_to_MUX_Product118_impl_0_parent_implementedSystem_port_1_cast <= SharedReg288_out;
SharedReg322_out_to_MUX_Product118_impl_0_parent_implementedSystem_port_2_cast <= SharedReg322_out;
   MUX_Product118_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg288_out_to_MUX_Product118_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg322_out_to_MUX_Product118_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product118_impl_0_out);

   Delay1No256_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product118_impl_0_out,
                 Y => Delay1No256_out);

SharedReg229_out_to_MUX_Product118_impl_1_parent_implementedSystem_port_1_cast <= SharedReg229_out;
SharedReg55_out_to_MUX_Product118_impl_1_parent_implementedSystem_port_2_cast <= SharedReg55_out;
   MUX_Product118_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg229_out_to_MUX_Product118_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg55_out_to_MUX_Product118_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product118_impl_1_out);

   Delay1No257_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product118_impl_1_out,
                 Y => Delay1No257_out);

Delay1No258_out_to_Product217_impl_parent_implementedSystem_port_0_cast <= Delay1No258_out;
Delay1No259_out_to_Product217_impl_parent_implementedSystem_port_1_cast <= Delay1No259_out;
   Product217_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product217_impl_out,
                 X => Delay1No258_out_to_Product217_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No259_out_to_Product217_impl_parent_implementedSystem_port_1_cast);

SharedReg289_out_to_MUX_Product217_impl_0_parent_implementedSystem_port_1_cast <= SharedReg289_out;
SharedReg323_out_to_MUX_Product217_impl_0_parent_implementedSystem_port_2_cast <= SharedReg323_out;
   MUX_Product217_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg289_out_to_MUX_Product217_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg323_out_to_MUX_Product217_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product217_impl_0_out);

   Delay1No258_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product217_impl_0_out,
                 Y => Delay1No258_out);

SharedReg228_out_to_MUX_Product217_impl_1_parent_implementedSystem_port_1_cast <= SharedReg228_out;
SharedReg53_out_to_MUX_Product217_impl_1_parent_implementedSystem_port_2_cast <= SharedReg53_out;
   MUX_Product217_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg228_out_to_MUX_Product217_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg53_out_to_MUX_Product217_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product217_impl_1_out);

   Delay1No259_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product217_impl_1_out,
                 Y => Delay1No259_out);

Delay1No260_out_to_Product317_impl_parent_implementedSystem_port_0_cast <= Delay1No260_out;
Delay1No261_out_to_Product317_impl_parent_implementedSystem_port_1_cast <= Delay1No261_out;
   Product317_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product317_impl_out,
                 X => Delay1No260_out_to_Product317_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No261_out_to_Product317_impl_parent_implementedSystem_port_1_cast);

SharedReg229_out_to_MUX_Product317_impl_0_parent_implementedSystem_port_1_cast <= SharedReg229_out;
SharedReg55_out_to_MUX_Product317_impl_0_parent_implementedSystem_port_2_cast <= SharedReg55_out;
   MUX_Product317_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg229_out_to_MUX_Product317_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg55_out_to_MUX_Product317_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product317_impl_0_out);

   Delay1No260_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product317_impl_0_out,
                 Y => Delay1No260_out);

SharedReg289_out_to_MUX_Product317_impl_1_parent_implementedSystem_port_1_cast <= SharedReg289_out;
SharedReg323_out_to_MUX_Product317_impl_1_parent_implementedSystem_port_2_cast <= SharedReg323_out;
   MUX_Product317_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg289_out_to_MUX_Product317_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg323_out_to_MUX_Product317_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product317_impl_1_out);

   Delay1No261_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product317_impl_1_out,
                 Y => Delay1No261_out);

Delay1No262_out_to_Subtract18_impl_parent_implementedSystem_port_0_cast <= Delay1No262_out;
Delay1No263_out_to_Subtract18_impl_parent_implementedSystem_port_1_cast <= Delay1No263_out;
   Subtract18_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract18_impl_out,
                 X => Delay1No262_out_to_Subtract18_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No263_out_to_Subtract18_impl_parent_implementedSystem_port_1_cast);

SharedReg155_out_to_MUX_Subtract18_impl_0_parent_implementedSystem_port_1_cast <= SharedReg155_out;
SharedReg161_out_to_MUX_Subtract18_impl_0_parent_implementedSystem_port_2_cast <= SharedReg161_out;
   MUX_Subtract18_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg155_out_to_MUX_Subtract18_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg161_out_to_MUX_Subtract18_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract18_impl_0_out);

   Delay1No262_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract18_impl_0_out,
                 Y => Delay1No262_out);

SharedReg158_out_to_MUX_Subtract18_impl_1_parent_implementedSystem_port_1_cast <= SharedReg158_out;
SharedReg164_out_to_MUX_Subtract18_impl_1_parent_implementedSystem_port_2_cast <= SharedReg164_out;
   MUX_Subtract18_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg158_out_to_MUX_Subtract18_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg164_out_to_MUX_Subtract18_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract18_impl_1_out);

   Delay1No263_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract18_impl_1_out,
                 Y => Delay1No263_out);

Delay1No264_out_to_Add61_impl_parent_implementedSystem_port_0_cast <= Delay1No264_out;
Delay1No265_out_to_Add61_impl_parent_implementedSystem_port_1_cast <= Delay1No265_out;
   Add61_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add61_impl_out,
                 X => Delay1No264_out_to_Add61_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No265_out_to_Add61_impl_parent_implementedSystem_port_1_cast);

SharedReg162_out_to_MUX_Add61_impl_0_parent_implementedSystem_port_1_cast <= SharedReg162_out;
SharedReg168_out_to_MUX_Add61_impl_0_parent_implementedSystem_port_2_cast <= SharedReg168_out;
   MUX_Add61_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg162_out_to_MUX_Add61_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg168_out_to_MUX_Add61_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add61_impl_0_out);

   Delay1No264_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add61_impl_0_out,
                 Y => Delay1No264_out);

SharedReg163_out_to_MUX_Add61_impl_1_parent_implementedSystem_port_1_cast <= SharedReg163_out;
SharedReg169_out_to_MUX_Add61_impl_1_parent_implementedSystem_port_2_cast <= SharedReg169_out;
   MUX_Add61_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg163_out_to_MUX_Add61_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg169_out_to_MUX_Add61_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add61_impl_1_out);

   Delay1No265_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add61_impl_1_out,
                 Y => Delay1No265_out);

Delay1No266_out_to_Product48_impl_parent_implementedSystem_port_0_cast <= Delay1No266_out;
Delay1No267_out_to_Product48_impl_parent_implementedSystem_port_1_cast <= Delay1No267_out;
   Product48_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product48_impl_out,
                 X => Delay1No266_out_to_Product48_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No267_out_to_Product48_impl_parent_implementedSystem_port_1_cast);

SharedReg292_out_to_MUX_Product48_impl_0_parent_implementedSystem_port_1_cast <= SharedReg292_out;
SharedReg328_out_to_MUX_Product48_impl_0_parent_implementedSystem_port_2_cast <= SharedReg328_out;
   MUX_Product48_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg292_out_to_MUX_Product48_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg328_out_to_MUX_Product48_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product48_impl_0_out);

   Delay1No266_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product48_impl_0_out,
                 Y => Delay1No266_out);

SharedReg35_out_to_MUX_Product48_impl_1_parent_implementedSystem_port_1_cast <= SharedReg35_out;
SharedReg57_out_to_MUX_Product48_impl_1_parent_implementedSystem_port_2_cast <= SharedReg57_out;
   MUX_Product48_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg35_out_to_MUX_Product48_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg57_out_to_MUX_Product48_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product48_impl_1_out);

   Delay1No267_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product48_impl_1_out,
                 Y => Delay1No267_out);

Delay1No268_out_to_Product120_impl_parent_implementedSystem_port_0_cast <= Delay1No268_out;
Delay1No269_out_to_Product120_impl_parent_implementedSystem_port_1_cast <= Delay1No269_out;
   Product120_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product120_impl_out,
                 X => Delay1No268_out_to_Product120_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No269_out_to_Product120_impl_parent_implementedSystem_port_1_cast);

SharedReg292_out_to_MUX_Product120_impl_0_parent_implementedSystem_port_1_cast <= SharedReg292_out;
SharedReg328_out_to_MUX_Product120_impl_0_parent_implementedSystem_port_2_cast <= SharedReg328_out;
   MUX_Product120_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg292_out_to_MUX_Product120_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg328_out_to_MUX_Product120_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product120_impl_0_out);

   Delay1No268_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product120_impl_0_out,
                 Y => Delay1No268_out);

SharedReg36_out_to_MUX_Product120_impl_1_parent_implementedSystem_port_1_cast <= SharedReg36_out;
SharedReg59_out_to_MUX_Product120_impl_1_parent_implementedSystem_port_2_cast <= SharedReg59_out;
   MUX_Product120_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg36_out_to_MUX_Product120_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg59_out_to_MUX_Product120_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product120_impl_1_out);

   Delay1No269_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product120_impl_1_out,
                 Y => Delay1No269_out);

Delay1No270_out_to_Product219_impl_parent_implementedSystem_port_0_cast <= Delay1No270_out;
Delay1No271_out_to_Product219_impl_parent_implementedSystem_port_1_cast <= Delay1No271_out;
   Product219_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product219_impl_out,
                 X => Delay1No270_out_to_Product219_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No271_out_to_Product219_impl_parent_implementedSystem_port_1_cast);

SharedReg293_out_to_MUX_Product219_impl_0_parent_implementedSystem_port_1_cast <= SharedReg293_out;
SharedReg329_out_to_MUX_Product219_impl_0_parent_implementedSystem_port_2_cast <= SharedReg329_out;
   MUX_Product219_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg293_out_to_MUX_Product219_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg329_out_to_MUX_Product219_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product219_impl_0_out);

   Delay1No270_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product219_impl_0_out,
                 Y => Delay1No270_out);

SharedReg35_out_to_MUX_Product219_impl_1_parent_implementedSystem_port_1_cast <= SharedReg35_out;
SharedReg57_out_to_MUX_Product219_impl_1_parent_implementedSystem_port_2_cast <= SharedReg57_out;
   MUX_Product219_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg35_out_to_MUX_Product219_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg57_out_to_MUX_Product219_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product219_impl_1_out);

   Delay1No271_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product219_impl_1_out,
                 Y => Delay1No271_out);

Delay1No272_out_to_Product319_impl_parent_implementedSystem_port_0_cast <= Delay1No272_out;
Delay1No273_out_to_Product319_impl_parent_implementedSystem_port_1_cast <= Delay1No273_out;
   Product319_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product319_impl_out,
                 X => Delay1No272_out_to_Product319_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No273_out_to_Product319_impl_parent_implementedSystem_port_1_cast);

SharedReg36_out_to_MUX_Product319_impl_0_parent_implementedSystem_port_1_cast <= SharedReg36_out;
SharedReg59_out_to_MUX_Product319_impl_0_parent_implementedSystem_port_2_cast <= SharedReg59_out;
   MUX_Product319_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg36_out_to_MUX_Product319_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg59_out_to_MUX_Product319_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product319_impl_0_out);

   Delay1No272_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product319_impl_0_out,
                 Y => Delay1No272_out);

SharedReg293_out_to_MUX_Product319_impl_1_parent_implementedSystem_port_1_cast <= SharedReg293_out;
SharedReg329_out_to_MUX_Product319_impl_1_parent_implementedSystem_port_2_cast <= SharedReg329_out;
   MUX_Product319_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg293_out_to_MUX_Product319_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg329_out_to_MUX_Product319_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product319_impl_1_out);

   Delay1No273_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product319_impl_1_out,
                 Y => Delay1No273_out);

Delay1No274_out_to_Subtract20_impl_parent_implementedSystem_port_0_cast <= Delay1No274_out;
Delay1No275_out_to_Subtract20_impl_parent_implementedSystem_port_1_cast <= Delay1No275_out;
   Subtract20_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract20_impl_out,
                 X => Delay1No274_out_to_Subtract20_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No275_out_to_Subtract20_impl_parent_implementedSystem_port_1_cast);

SharedReg161_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_1_cast <= SharedReg161_out;
SharedReg167_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_2_cast <= SharedReg167_out;
   MUX_Subtract20_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg161_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg167_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract20_impl_0_out);

   Delay1No274_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract20_impl_0_out,
                 Y => Delay1No274_out);

SharedReg164_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_1_cast <= SharedReg164_out;
SharedReg170_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_2_cast <= SharedReg170_out;
   MUX_Subtract20_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg164_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg170_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract20_impl_1_out);

   Delay1No275_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract20_impl_1_out,
                 Y => Delay1No275_out);

Delay1No276_out_to_Add63_impl_parent_implementedSystem_port_0_cast <= Delay1No276_out;
Delay1No277_out_to_Add63_impl_parent_implementedSystem_port_1_cast <= Delay1No277_out;
   Add63_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add63_impl_out,
                 X => Delay1No276_out_to_Add63_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No277_out_to_Add63_impl_parent_implementedSystem_port_1_cast);

SharedReg168_out_to_MUX_Add63_impl_0_parent_implementedSystem_port_1_cast <= SharedReg168_out;
SharedReg174_out_to_MUX_Add63_impl_0_parent_implementedSystem_port_2_cast <= SharedReg174_out;
   MUX_Add63_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg168_out_to_MUX_Add63_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg174_out_to_MUX_Add63_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add63_impl_0_out);

   Delay1No276_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add63_impl_0_out,
                 Y => Delay1No276_out);

SharedReg169_out_to_MUX_Add63_impl_1_parent_implementedSystem_port_1_cast <= SharedReg169_out;
SharedReg175_out_to_MUX_Add63_impl_1_parent_implementedSystem_port_2_cast <= SharedReg175_out;
   MUX_Add63_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg169_out_to_MUX_Add63_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg175_out_to_MUX_Add63_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add63_impl_1_out);

   Delay1No277_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add63_impl_1_out,
                 Y => Delay1No277_out);

Delay1No278_out_to_Product50_impl_parent_implementedSystem_port_0_cast <= Delay1No278_out;
Delay1No279_out_to_Product50_impl_parent_implementedSystem_port_1_cast <= Delay1No279_out;
   Product50_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product50_impl_out,
                 X => Delay1No278_out_to_Product50_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No279_out_to_Product50_impl_parent_implementedSystem_port_1_cast);

SharedReg296_out_to_MUX_Product50_impl_0_parent_implementedSystem_port_1_cast <= SharedReg296_out;
SharedReg324_out_to_MUX_Product50_impl_0_parent_implementedSystem_port_2_cast <= SharedReg324_out;
   MUX_Product50_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg296_out_to_MUX_Product50_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg324_out_to_MUX_Product50_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product50_impl_0_out);

   Delay1No278_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product50_impl_0_out,
                 Y => Delay1No278_out);

SharedReg254_out_to_MUX_Product50_impl_1_parent_implementedSystem_port_1_cast <= SharedReg254_out;
SharedReg71_out_to_MUX_Product50_impl_1_parent_implementedSystem_port_2_cast <= SharedReg71_out;
   MUX_Product50_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg254_out_to_MUX_Product50_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg71_out_to_MUX_Product50_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product50_impl_1_out);

   Delay1No279_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product50_impl_1_out,
                 Y => Delay1No279_out);

Delay1No280_out_to_Product122_impl_parent_implementedSystem_port_0_cast <= Delay1No280_out;
Delay1No281_out_to_Product122_impl_parent_implementedSystem_port_1_cast <= Delay1No281_out;
   Product122_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product122_impl_out,
                 X => Delay1No280_out_to_Product122_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No281_out_to_Product122_impl_parent_implementedSystem_port_1_cast);

SharedReg296_out_to_MUX_Product122_impl_0_parent_implementedSystem_port_1_cast <= SharedReg296_out;
SharedReg324_out_to_MUX_Product122_impl_0_parent_implementedSystem_port_2_cast <= SharedReg324_out;
   MUX_Product122_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg296_out_to_MUX_Product122_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg324_out_to_MUX_Product122_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product122_impl_0_out);

   Delay1No280_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product122_impl_0_out,
                 Y => Delay1No280_out);

SharedReg255_out_to_MUX_Product122_impl_1_parent_implementedSystem_port_1_cast <= SharedReg255_out;
SharedReg72_out_to_MUX_Product122_impl_1_parent_implementedSystem_port_2_cast <= SharedReg72_out;
   MUX_Product122_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg255_out_to_MUX_Product122_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg72_out_to_MUX_Product122_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product122_impl_1_out);

   Delay1No281_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product122_impl_1_out,
                 Y => Delay1No281_out);

Delay1No282_out_to_Product221_impl_parent_implementedSystem_port_0_cast <= Delay1No282_out;
Delay1No283_out_to_Product221_impl_parent_implementedSystem_port_1_cast <= Delay1No283_out;
   Product221_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product221_impl_out,
                 X => Delay1No282_out_to_Product221_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No283_out_to_Product221_impl_parent_implementedSystem_port_1_cast);

SharedReg297_out_to_MUX_Product221_impl_0_parent_implementedSystem_port_1_cast <= SharedReg297_out;
SharedReg325_out_to_MUX_Product221_impl_0_parent_implementedSystem_port_2_cast <= SharedReg325_out;
   MUX_Product221_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg297_out_to_MUX_Product221_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg325_out_to_MUX_Product221_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product221_impl_0_out);

   Delay1No282_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product221_impl_0_out,
                 Y => Delay1No282_out);

SharedReg254_out_to_MUX_Product221_impl_1_parent_implementedSystem_port_1_cast <= SharedReg254_out;
SharedReg71_out_to_MUX_Product221_impl_1_parent_implementedSystem_port_2_cast <= SharedReg71_out;
   MUX_Product221_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg254_out_to_MUX_Product221_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg71_out_to_MUX_Product221_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product221_impl_1_out);

   Delay1No283_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product221_impl_1_out,
                 Y => Delay1No283_out);

Delay1No284_out_to_Product321_impl_parent_implementedSystem_port_0_cast <= Delay1No284_out;
Delay1No285_out_to_Product321_impl_parent_implementedSystem_port_1_cast <= Delay1No285_out;
   Product321_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product321_impl_out,
                 X => Delay1No284_out_to_Product321_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No285_out_to_Product321_impl_parent_implementedSystem_port_1_cast);

SharedReg255_out_to_MUX_Product321_impl_0_parent_implementedSystem_port_1_cast <= SharedReg255_out;
SharedReg72_out_to_MUX_Product321_impl_0_parent_implementedSystem_port_2_cast <= SharedReg72_out;
   MUX_Product321_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg255_out_to_MUX_Product321_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg72_out_to_MUX_Product321_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product321_impl_0_out);

   Delay1No284_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_impl_0_out,
                 Y => Delay1No284_out);

SharedReg297_out_to_MUX_Product321_impl_1_parent_implementedSystem_port_1_cast <= SharedReg297_out;
SharedReg325_out_to_MUX_Product321_impl_1_parent_implementedSystem_port_2_cast <= SharedReg325_out;
   MUX_Product321_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg297_out_to_MUX_Product321_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg325_out_to_MUX_Product321_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product321_impl_1_out);

   Delay1No285_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_impl_1_out,
                 Y => Delay1No285_out);

Delay1No286_out_to_Subtract22_impl_parent_implementedSystem_port_0_cast <= Delay1No286_out;
Delay1No287_out_to_Subtract22_impl_parent_implementedSystem_port_1_cast <= Delay1No287_out;
   Subtract22_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract22_impl_out,
                 X => Delay1No286_out_to_Subtract22_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No287_out_to_Subtract22_impl_parent_implementedSystem_port_1_cast);

SharedReg167_out_to_MUX_Subtract22_impl_0_parent_implementedSystem_port_1_cast <= SharedReg167_out;
SharedReg173_out_to_MUX_Subtract22_impl_0_parent_implementedSystem_port_2_cast <= SharedReg173_out;
   MUX_Subtract22_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg167_out_to_MUX_Subtract22_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg173_out_to_MUX_Subtract22_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract22_impl_0_out);

   Delay1No286_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract22_impl_0_out,
                 Y => Delay1No286_out);

SharedReg170_out_to_MUX_Subtract22_impl_1_parent_implementedSystem_port_1_cast <= SharedReg170_out;
SharedReg176_out_to_MUX_Subtract22_impl_1_parent_implementedSystem_port_2_cast <= SharedReg176_out;
   MUX_Subtract22_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg170_out_to_MUX_Subtract22_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg176_out_to_MUX_Subtract22_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract22_impl_1_out);

   Delay1No287_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract22_impl_1_out,
                 Y => Delay1No287_out);

Delay1No288_out_to_Add65_impl_parent_implementedSystem_port_0_cast <= Delay1No288_out;
Delay1No289_out_to_Add65_impl_parent_implementedSystem_port_1_cast <= Delay1No289_out;
   Add65_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add65_impl_out,
                 X => Delay1No288_out_to_Add65_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No289_out_to_Add65_impl_parent_implementedSystem_port_1_cast);

SharedReg174_out_to_MUX_Add65_impl_0_parent_implementedSystem_port_1_cast <= SharedReg174_out;
SharedReg180_out_to_MUX_Add65_impl_0_parent_implementedSystem_port_2_cast <= SharedReg180_out;
   MUX_Add65_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg174_out_to_MUX_Add65_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg180_out_to_MUX_Add65_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add65_impl_0_out);

   Delay1No288_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add65_impl_0_out,
                 Y => Delay1No288_out);

SharedReg175_out_to_MUX_Add65_impl_1_parent_implementedSystem_port_1_cast <= SharedReg175_out;
SharedReg181_out_to_MUX_Add65_impl_1_parent_implementedSystem_port_2_cast <= SharedReg181_out;
   MUX_Add65_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg175_out_to_MUX_Add65_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg181_out_to_MUX_Add65_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add65_impl_1_out);

   Delay1No289_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add65_impl_1_out,
                 Y => Delay1No289_out);

Delay1No290_out_to_Product52_impl_parent_implementedSystem_port_0_cast <= Delay1No290_out;
Delay1No291_out_to_Product52_impl_parent_implementedSystem_port_1_cast <= Delay1No291_out;
   Product52_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product52_impl_out,
                 X => Delay1No290_out_to_Product52_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No291_out_to_Product52_impl_parent_implementedSystem_port_1_cast);

SharedReg268_out_to_MUX_Product52_impl_0_parent_implementedSystem_port_1_cast <= SharedReg268_out;
SharedReg326_out_to_MUX_Product52_impl_0_parent_implementedSystem_port_2_cast <= SharedReg326_out;
   MUX_Product52_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg268_out_to_MUX_Product52_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg326_out_to_MUX_Product52_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product52_impl_0_out);

   Delay1No290_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product52_impl_0_out,
                 Y => Delay1No290_out);

SharedReg223_out_to_MUX_Product52_impl_1_parent_implementedSystem_port_1_cast <= SharedReg223_out;
SharedReg227_out_to_MUX_Product52_impl_1_parent_implementedSystem_port_2_cast <= SharedReg227_out;
   MUX_Product52_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg223_out_to_MUX_Product52_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg227_out_to_MUX_Product52_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product52_impl_1_out);

   Delay1No291_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product52_impl_1_out,
                 Y => Delay1No291_out);

Delay1No292_out_to_Product124_impl_parent_implementedSystem_port_0_cast <= Delay1No292_out;
Delay1No293_out_to_Product124_impl_parent_implementedSystem_port_1_cast <= Delay1No293_out;
   Product124_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product124_impl_out,
                 X => Delay1No292_out_to_Product124_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No293_out_to_Product124_impl_parent_implementedSystem_port_1_cast);

SharedReg268_out_to_MUX_Product124_impl_0_parent_implementedSystem_port_1_cast <= SharedReg268_out;
SharedReg326_out_to_MUX_Product124_impl_0_parent_implementedSystem_port_2_cast <= SharedReg326_out;
   MUX_Product124_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg268_out_to_MUX_Product124_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg326_out_to_MUX_Product124_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product124_impl_0_out);

   Delay1No292_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product124_impl_0_out,
                 Y => Delay1No292_out);

SharedReg225_out_to_MUX_Product124_impl_1_parent_implementedSystem_port_1_cast <= SharedReg225_out;
SharedReg228_out_to_MUX_Product124_impl_1_parent_implementedSystem_port_2_cast <= SharedReg228_out;
   MUX_Product124_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg225_out_to_MUX_Product124_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg228_out_to_MUX_Product124_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product124_impl_1_out);

   Delay1No293_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product124_impl_1_out,
                 Y => Delay1No293_out);

Delay1No294_out_to_Product223_impl_parent_implementedSystem_port_0_cast <= Delay1No294_out;
Delay1No295_out_to_Product223_impl_parent_implementedSystem_port_1_cast <= Delay1No295_out;
   Product223_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product223_impl_out,
                 X => Delay1No294_out_to_Product223_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No295_out_to_Product223_impl_parent_implementedSystem_port_1_cast);

SharedReg269_out_to_MUX_Product223_impl_0_parent_implementedSystem_port_1_cast <= SharedReg269_out;
SharedReg327_out_to_MUX_Product223_impl_0_parent_implementedSystem_port_2_cast <= SharedReg327_out;
   MUX_Product223_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg269_out_to_MUX_Product223_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg327_out_to_MUX_Product223_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product223_impl_0_out);

   Delay1No294_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product223_impl_0_out,
                 Y => Delay1No294_out);

SharedReg223_out_to_MUX_Product223_impl_1_parent_implementedSystem_port_1_cast <= SharedReg223_out;
SharedReg227_out_to_MUX_Product223_impl_1_parent_implementedSystem_port_2_cast <= SharedReg227_out;
   MUX_Product223_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg223_out_to_MUX_Product223_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg227_out_to_MUX_Product223_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product223_impl_1_out);

   Delay1No295_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product223_impl_1_out,
                 Y => Delay1No295_out);

Delay1No296_out_to_Product323_impl_parent_implementedSystem_port_0_cast <= Delay1No296_out;
Delay1No297_out_to_Product323_impl_parent_implementedSystem_port_1_cast <= Delay1No297_out;
   Product323_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product323_impl_out,
                 X => Delay1No296_out_to_Product323_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No297_out_to_Product323_impl_parent_implementedSystem_port_1_cast);

SharedReg225_out_to_MUX_Product323_impl_0_parent_implementedSystem_port_1_cast <= SharedReg225_out;
SharedReg228_out_to_MUX_Product323_impl_0_parent_implementedSystem_port_2_cast <= SharedReg228_out;
   MUX_Product323_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg225_out_to_MUX_Product323_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg228_out_to_MUX_Product323_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product323_impl_0_out);

   Delay1No296_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product323_impl_0_out,
                 Y => Delay1No296_out);

SharedReg269_out_to_MUX_Product323_impl_1_parent_implementedSystem_port_1_cast <= SharedReg269_out;
SharedReg327_out_to_MUX_Product323_impl_1_parent_implementedSystem_port_2_cast <= SharedReg327_out;
   MUX_Product323_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg269_out_to_MUX_Product323_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg327_out_to_MUX_Product323_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product323_impl_1_out);

   Delay1No297_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product323_impl_1_out,
                 Y => Delay1No297_out);

Delay1No298_out_to_Subtract24_impl_parent_implementedSystem_port_0_cast <= Delay1No298_out;
Delay1No299_out_to_Subtract24_impl_parent_implementedSystem_port_1_cast <= Delay1No299_out;
   Subtract24_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract24_impl_out,
                 X => Delay1No298_out_to_Subtract24_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No299_out_to_Subtract24_impl_parent_implementedSystem_port_1_cast);

SharedReg173_out_to_MUX_Subtract24_impl_0_parent_implementedSystem_port_1_cast <= SharedReg173_out;
SharedReg179_out_to_MUX_Subtract24_impl_0_parent_implementedSystem_port_2_cast <= SharedReg179_out;
   MUX_Subtract24_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg173_out_to_MUX_Subtract24_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg179_out_to_MUX_Subtract24_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract24_impl_0_out);

   Delay1No298_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract24_impl_0_out,
                 Y => Delay1No298_out);

SharedReg176_out_to_MUX_Subtract24_impl_1_parent_implementedSystem_port_1_cast <= SharedReg176_out;
SharedReg182_out_to_MUX_Subtract24_impl_1_parent_implementedSystem_port_2_cast <= SharedReg182_out;
   MUX_Subtract24_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg176_out_to_MUX_Subtract24_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg182_out_to_MUX_Subtract24_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract24_impl_1_out);

   Delay1No299_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract24_impl_1_out,
                 Y => Delay1No299_out);

Delay1No300_out_to_Add66_impl_parent_implementedSystem_port_0_cast <= Delay1No300_out;
Delay1No301_out_to_Add66_impl_parent_implementedSystem_port_1_cast <= Delay1No301_out;
   Add66_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add66_impl_out,
                 X => Delay1No300_out_to_Add66_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No301_out_to_Add66_impl_parent_implementedSystem_port_1_cast);

SharedReg180_out_to_MUX_Add66_impl_0_parent_implementedSystem_port_1_cast <= SharedReg180_out;
SharedReg186_out_to_MUX_Add66_impl_0_parent_implementedSystem_port_2_cast <= SharedReg186_out;
   MUX_Add66_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg180_out_to_MUX_Add66_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg186_out_to_MUX_Add66_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add66_impl_0_out);

   Delay1No300_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add66_impl_0_out,
                 Y => Delay1No300_out);

SharedReg181_out_to_MUX_Add66_impl_1_parent_implementedSystem_port_1_cast <= SharedReg181_out;
SharedReg187_out_to_MUX_Add66_impl_1_parent_implementedSystem_port_2_cast <= SharedReg187_out;
   MUX_Add66_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg181_out_to_MUX_Add66_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg187_out_to_MUX_Add66_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add66_impl_1_out);

   Delay1No301_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add66_impl_1_out,
                 Y => Delay1No301_out);

Delay1No302_out_to_Product53_impl_parent_implementedSystem_port_0_cast <= Delay1No302_out;
Delay1No303_out_to_Product53_impl_parent_implementedSystem_port_1_cast <= Delay1No303_out;
   Product53_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product53_impl_out,
                 X => Delay1No302_out_to_Product53_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No303_out_to_Product53_impl_parent_implementedSystem_port_1_cast);

SharedReg302_out_to_MUX_Product53_impl_0_parent_implementedSystem_port_1_cast <= SharedReg302_out;
SharedReg312_out_to_MUX_Product53_impl_0_parent_implementedSystem_port_2_cast <= SharedReg312_out;
   MUX_Product53_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg302_out_to_MUX_Product53_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg312_out_to_MUX_Product53_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product53_impl_0_out);

   Delay1No302_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product53_impl_0_out,
                 Y => Delay1No302_out);

SharedReg68_out_to_MUX_Product53_impl_1_parent_implementedSystem_port_1_cast <= SharedReg68_out;
SharedReg235_out_to_MUX_Product53_impl_1_parent_implementedSystem_port_2_cast <= SharedReg235_out;
   MUX_Product53_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg68_out_to_MUX_Product53_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg235_out_to_MUX_Product53_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product53_impl_1_out);

   Delay1No303_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product53_impl_1_out,
                 Y => Delay1No303_out);

Delay1No304_out_to_Product125_impl_parent_implementedSystem_port_0_cast <= Delay1No304_out;
Delay1No305_out_to_Product125_impl_parent_implementedSystem_port_1_cast <= Delay1No305_out;
   Product125_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product125_impl_out,
                 X => Delay1No304_out_to_Product125_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No305_out_to_Product125_impl_parent_implementedSystem_port_1_cast);

SharedReg302_out_to_MUX_Product125_impl_0_parent_implementedSystem_port_1_cast <= SharedReg302_out;
SharedReg312_out_to_MUX_Product125_impl_0_parent_implementedSystem_port_2_cast <= SharedReg312_out;
   MUX_Product125_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg302_out_to_MUX_Product125_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg312_out_to_MUX_Product125_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product125_impl_0_out);

   Delay1No304_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product125_impl_0_out,
                 Y => Delay1No304_out);

SharedReg69_out_to_MUX_Product125_impl_1_parent_implementedSystem_port_1_cast <= SharedReg69_out;
SharedReg237_out_to_MUX_Product125_impl_1_parent_implementedSystem_port_2_cast <= SharedReg237_out;
   MUX_Product125_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg69_out_to_MUX_Product125_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg237_out_to_MUX_Product125_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product125_impl_1_out);

   Delay1No305_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product125_impl_1_out,
                 Y => Delay1No305_out);

Delay1No306_out_to_Product224_impl_parent_implementedSystem_port_0_cast <= Delay1No306_out;
Delay1No307_out_to_Product224_impl_parent_implementedSystem_port_1_cast <= Delay1No307_out;
   Product224_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product224_impl_out,
                 X => Delay1No306_out_to_Product224_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No307_out_to_Product224_impl_parent_implementedSystem_port_1_cast);

SharedReg303_out_to_MUX_Product224_impl_0_parent_implementedSystem_port_1_cast <= SharedReg303_out;
SharedReg313_out_to_MUX_Product224_impl_0_parent_implementedSystem_port_2_cast <= SharedReg313_out;
   MUX_Product224_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg303_out_to_MUX_Product224_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg313_out_to_MUX_Product224_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product224_impl_0_out);

   Delay1No306_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product224_impl_0_out,
                 Y => Delay1No306_out);

SharedReg68_out_to_MUX_Product224_impl_1_parent_implementedSystem_port_1_cast <= SharedReg68_out;
SharedReg235_out_to_MUX_Product224_impl_1_parent_implementedSystem_port_2_cast <= SharedReg235_out;
   MUX_Product224_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg68_out_to_MUX_Product224_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg235_out_to_MUX_Product224_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product224_impl_1_out);

   Delay1No307_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product224_impl_1_out,
                 Y => Delay1No307_out);

Delay1No308_out_to_Product324_impl_parent_implementedSystem_port_0_cast <= Delay1No308_out;
Delay1No309_out_to_Product324_impl_parent_implementedSystem_port_1_cast <= Delay1No309_out;
   Product324_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product324_impl_out,
                 X => Delay1No308_out_to_Product324_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No309_out_to_Product324_impl_parent_implementedSystem_port_1_cast);

SharedReg69_out_to_MUX_Product324_impl_0_parent_implementedSystem_port_1_cast <= SharedReg69_out;
SharedReg237_out_to_MUX_Product324_impl_0_parent_implementedSystem_port_2_cast <= SharedReg237_out;
   MUX_Product324_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg69_out_to_MUX_Product324_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg237_out_to_MUX_Product324_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product324_impl_0_out);

   Delay1No308_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product324_impl_0_out,
                 Y => Delay1No308_out);

SharedReg303_out_to_MUX_Product324_impl_1_parent_implementedSystem_port_1_cast <= SharedReg303_out;
SharedReg313_out_to_MUX_Product324_impl_1_parent_implementedSystem_port_2_cast <= SharedReg313_out;
   MUX_Product324_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg303_out_to_MUX_Product324_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg313_out_to_MUX_Product324_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product324_impl_1_out);

   Delay1No309_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product324_impl_1_out,
                 Y => Delay1No309_out);

Delay1No310_out_to_Subtract25_impl_parent_implementedSystem_port_0_cast <= Delay1No310_out;
Delay1No311_out_to_Subtract25_impl_parent_implementedSystem_port_1_cast <= Delay1No311_out;
   Subtract25_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract25_impl_out,
                 X => Delay1No310_out_to_Subtract25_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No311_out_to_Subtract25_impl_parent_implementedSystem_port_1_cast);

SharedReg179_out_to_MUX_Subtract25_impl_0_parent_implementedSystem_port_1_cast <= SharedReg179_out;
SharedReg185_out_to_MUX_Subtract25_impl_0_parent_implementedSystem_port_2_cast <= SharedReg185_out;
   MUX_Subtract25_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg179_out_to_MUX_Subtract25_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg185_out_to_MUX_Subtract25_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract25_impl_0_out);

   Delay1No310_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract25_impl_0_out,
                 Y => Delay1No310_out);

SharedReg182_out_to_MUX_Subtract25_impl_1_parent_implementedSystem_port_1_cast <= SharedReg182_out;
SharedReg188_out_to_MUX_Subtract25_impl_1_parent_implementedSystem_port_2_cast <= SharedReg188_out;
   MUX_Subtract25_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg182_out_to_MUX_Subtract25_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg188_out_to_MUX_Subtract25_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract25_impl_1_out);

   Delay1No311_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract25_impl_1_out,
                 Y => Delay1No311_out);

Delay1No312_out_to_Add67_impl_parent_implementedSystem_port_0_cast <= Delay1No312_out;
Delay1No313_out_to_Add67_impl_parent_implementedSystem_port_1_cast <= Delay1No313_out;
   Add67_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add67_impl_out,
                 X => Delay1No312_out_to_Add67_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No313_out_to_Add67_impl_parent_implementedSystem_port_1_cast);

SharedReg186_out_to_MUX_Add67_impl_0_parent_implementedSystem_port_1_cast <= SharedReg186_out;
SharedReg192_out_to_MUX_Add67_impl_0_parent_implementedSystem_port_2_cast <= SharedReg192_out;
   MUX_Add67_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg186_out_to_MUX_Add67_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg192_out_to_MUX_Add67_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add67_impl_0_out);

   Delay1No312_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add67_impl_0_out,
                 Y => Delay1No312_out);

SharedReg187_out_to_MUX_Add67_impl_1_parent_implementedSystem_port_1_cast <= SharedReg187_out;
SharedReg193_out_to_MUX_Add67_impl_1_parent_implementedSystem_port_2_cast <= SharedReg193_out;
   MUX_Add67_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg187_out_to_MUX_Add67_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg193_out_to_MUX_Add67_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add67_impl_1_out);

   Delay1No313_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add67_impl_1_out,
                 Y => Delay1No313_out);

Delay1No314_out_to_Product54_impl_parent_implementedSystem_port_0_cast <= Delay1No314_out;
Delay1No315_out_to_Product54_impl_parent_implementedSystem_port_1_cast <= Delay1No315_out;
   Product54_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product54_impl_out,
                 X => Delay1No314_out_to_Product54_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No315_out_to_Product54_impl_parent_implementedSystem_port_1_cast);

SharedReg304_out_to_MUX_Product54_impl_0_parent_implementedSystem_port_1_cast <= SharedReg304_out;
SharedReg332_out_to_MUX_Product54_impl_0_parent_implementedSystem_port_2_cast <= SharedReg332_out;
   MUX_Product54_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg304_out_to_MUX_Product54_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg332_out_to_MUX_Product54_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product54_impl_0_out);

   Delay1No314_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product54_impl_0_out,
                 Y => Delay1No314_out);

SharedReg230_out_to_MUX_Product54_impl_1_parent_implementedSystem_port_1_cast <= SharedReg230_out;
SharedReg241_out_to_MUX_Product54_impl_1_parent_implementedSystem_port_2_cast <= SharedReg241_out;
   MUX_Product54_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg230_out_to_MUX_Product54_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg241_out_to_MUX_Product54_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product54_impl_1_out);

   Delay1No315_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product54_impl_1_out,
                 Y => Delay1No315_out);

Delay1No316_out_to_Product126_impl_parent_implementedSystem_port_0_cast <= Delay1No316_out;
Delay1No317_out_to_Product126_impl_parent_implementedSystem_port_1_cast <= Delay1No317_out;
   Product126_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product126_impl_out,
                 X => Delay1No316_out_to_Product126_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No317_out_to_Product126_impl_parent_implementedSystem_port_1_cast);

SharedReg304_out_to_MUX_Product126_impl_0_parent_implementedSystem_port_1_cast <= SharedReg304_out;
SharedReg332_out_to_MUX_Product126_impl_0_parent_implementedSystem_port_2_cast <= SharedReg332_out;
   MUX_Product126_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg304_out_to_MUX_Product126_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg332_out_to_MUX_Product126_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product126_impl_0_out);

   Delay1No316_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product126_impl_0_out,
                 Y => Delay1No316_out);

SharedReg231_out_to_MUX_Product126_impl_1_parent_implementedSystem_port_1_cast <= SharedReg231_out;
SharedReg243_out_to_MUX_Product126_impl_1_parent_implementedSystem_port_2_cast <= SharedReg243_out;
   MUX_Product126_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg231_out_to_MUX_Product126_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg243_out_to_MUX_Product126_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product126_impl_1_out);

   Delay1No317_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product126_impl_1_out,
                 Y => Delay1No317_out);

Delay1No318_out_to_Product225_impl_parent_implementedSystem_port_0_cast <= Delay1No318_out;
Delay1No319_out_to_Product225_impl_parent_implementedSystem_port_1_cast <= Delay1No319_out;
   Product225_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product225_impl_out,
                 X => Delay1No318_out_to_Product225_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No319_out_to_Product225_impl_parent_implementedSystem_port_1_cast);

SharedReg305_out_to_MUX_Product225_impl_0_parent_implementedSystem_port_1_cast <= SharedReg305_out;
SharedReg333_out_to_MUX_Product225_impl_0_parent_implementedSystem_port_2_cast <= SharedReg333_out;
   MUX_Product225_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg305_out_to_MUX_Product225_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg333_out_to_MUX_Product225_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product225_impl_0_out);

   Delay1No318_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product225_impl_0_out,
                 Y => Delay1No318_out);

SharedReg230_out_to_MUX_Product225_impl_1_parent_implementedSystem_port_1_cast <= SharedReg230_out;
SharedReg241_out_to_MUX_Product225_impl_1_parent_implementedSystem_port_2_cast <= SharedReg241_out;
   MUX_Product225_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg230_out_to_MUX_Product225_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg241_out_to_MUX_Product225_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product225_impl_1_out);

   Delay1No319_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product225_impl_1_out,
                 Y => Delay1No319_out);

Delay1No320_out_to_Product325_impl_parent_implementedSystem_port_0_cast <= Delay1No320_out;
Delay1No321_out_to_Product325_impl_parent_implementedSystem_port_1_cast <= Delay1No321_out;
   Product325_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product325_impl_out,
                 X => Delay1No320_out_to_Product325_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No321_out_to_Product325_impl_parent_implementedSystem_port_1_cast);

SharedReg231_out_to_MUX_Product325_impl_0_parent_implementedSystem_port_1_cast <= SharedReg231_out;
SharedReg243_out_to_MUX_Product325_impl_0_parent_implementedSystem_port_2_cast <= SharedReg243_out;
   MUX_Product325_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg231_out_to_MUX_Product325_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg243_out_to_MUX_Product325_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product325_impl_0_out);

   Delay1No320_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product325_impl_0_out,
                 Y => Delay1No320_out);

SharedReg305_out_to_MUX_Product325_impl_1_parent_implementedSystem_port_1_cast <= SharedReg305_out;
SharedReg333_out_to_MUX_Product325_impl_1_parent_implementedSystem_port_2_cast <= SharedReg333_out;
   MUX_Product325_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg305_out_to_MUX_Product325_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg333_out_to_MUX_Product325_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product325_impl_1_out);

   Delay1No321_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product325_impl_1_out,
                 Y => Delay1No321_out);

Delay1No322_out_to_Subtract26_impl_parent_implementedSystem_port_0_cast <= Delay1No322_out;
Delay1No323_out_to_Subtract26_impl_parent_implementedSystem_port_1_cast <= Delay1No323_out;
   Subtract26_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract26_impl_out,
                 X => Delay1No322_out_to_Subtract26_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No323_out_to_Subtract26_impl_parent_implementedSystem_port_1_cast);

SharedReg185_out_to_MUX_Subtract26_impl_0_parent_implementedSystem_port_1_cast <= SharedReg185_out;
SharedReg191_out_to_MUX_Subtract26_impl_0_parent_implementedSystem_port_2_cast <= SharedReg191_out;
   MUX_Subtract26_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg185_out_to_MUX_Subtract26_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg191_out_to_MUX_Subtract26_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract26_impl_0_out);

   Delay1No322_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract26_impl_0_out,
                 Y => Delay1No322_out);

SharedReg188_out_to_MUX_Subtract26_impl_1_parent_implementedSystem_port_1_cast <= SharedReg188_out;
SharedReg194_out_to_MUX_Subtract26_impl_1_parent_implementedSystem_port_2_cast <= SharedReg194_out;
   MUX_Subtract26_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg188_out_to_MUX_Subtract26_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg194_out_to_MUX_Subtract26_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract26_impl_1_out);

   Delay1No323_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract26_impl_1_out,
                 Y => Delay1No323_out);

Delay1No324_out_to_Add68_impl_parent_implementedSystem_port_0_cast <= Delay1No324_out;
Delay1No325_out_to_Add68_impl_parent_implementedSystem_port_1_cast <= Delay1No325_out;
   Add68_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add68_impl_out,
                 X => Delay1No324_out_to_Add68_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No325_out_to_Add68_impl_parent_implementedSystem_port_1_cast);

SharedReg192_out_to_MUX_Add68_impl_0_parent_implementedSystem_port_1_cast <= SharedReg192_out;
SharedReg125_out_to_MUX_Add68_impl_0_parent_implementedSystem_port_2_cast <= SharedReg125_out;
   MUX_Add68_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg192_out_to_MUX_Add68_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg125_out_to_MUX_Add68_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add68_impl_0_out);

   Delay1No324_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add68_impl_0_out,
                 Y => Delay1No324_out);

SharedReg193_out_to_MUX_Add68_impl_1_parent_implementedSystem_port_1_cast <= SharedReg193_out;
SharedReg126_out_to_MUX_Add68_impl_1_parent_implementedSystem_port_2_cast <= SharedReg126_out;
   MUX_Add68_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg193_out_to_MUX_Add68_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg126_out_to_MUX_Add68_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add68_impl_1_out);

   Delay1No325_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add68_impl_1_out,
                 Y => Delay1No325_out);

Delay1No326_out_to_Product55_impl_parent_implementedSystem_port_0_cast <= Delay1No326_out;
Delay1No327_out_to_Product55_impl_parent_implementedSystem_port_1_cast <= Delay1No327_out;
   Product55_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product55_impl_out,
                 X => Delay1No326_out_to_Product55_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No327_out_to_Product55_impl_parent_implementedSystem_port_1_cast);

SharedReg298_out_to_MUX_Product55_impl_0_parent_implementedSystem_port_1_cast <= SharedReg298_out;
SharedReg330_out_to_MUX_Product55_impl_0_parent_implementedSystem_port_2_cast <= SharedReg330_out;
   MUX_Product55_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg298_out_to_MUX_Product55_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg330_out_to_MUX_Product55_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product55_impl_0_out);

   Delay1No326_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product55_impl_0_out,
                 Y => Delay1No326_out);

SharedReg232_out_to_MUX_Product55_impl_1_parent_implementedSystem_port_1_cast <= SharedReg232_out;
SharedReg233_out_to_MUX_Product55_impl_1_parent_implementedSystem_port_2_cast <= SharedReg233_out;
   MUX_Product55_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg232_out_to_MUX_Product55_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg233_out_to_MUX_Product55_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product55_impl_1_out);

   Delay1No327_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product55_impl_1_out,
                 Y => Delay1No327_out);

Delay1No328_out_to_Product127_impl_parent_implementedSystem_port_0_cast <= Delay1No328_out;
Delay1No329_out_to_Product127_impl_parent_implementedSystem_port_1_cast <= Delay1No329_out;
   Product127_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product127_impl_out,
                 X => Delay1No328_out_to_Product127_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No329_out_to_Product127_impl_parent_implementedSystem_port_1_cast);

SharedReg298_out_to_MUX_Product127_impl_0_parent_implementedSystem_port_1_cast <= SharedReg298_out;
SharedReg330_out_to_MUX_Product127_impl_0_parent_implementedSystem_port_2_cast <= SharedReg330_out;
   MUX_Product127_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg298_out_to_MUX_Product127_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg330_out_to_MUX_Product127_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product127_impl_0_out);

   Delay1No328_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product127_impl_0_out,
                 Y => Delay1No328_out);

SharedReg233_out_to_MUX_Product127_impl_1_parent_implementedSystem_port_1_cast <= SharedReg233_out;
SharedReg234_out_to_MUX_Product127_impl_1_parent_implementedSystem_port_2_cast <= SharedReg234_out;
   MUX_Product127_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg233_out_to_MUX_Product127_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg234_out_to_MUX_Product127_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product127_impl_1_out);

   Delay1No329_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product127_impl_1_out,
                 Y => Delay1No329_out);

Delay1No330_out_to_Product226_impl_parent_implementedSystem_port_0_cast <= Delay1No330_out;
Delay1No331_out_to_Product226_impl_parent_implementedSystem_port_1_cast <= Delay1No331_out;
   Product226_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product226_impl_out,
                 X => Delay1No330_out_to_Product226_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No331_out_to_Product226_impl_parent_implementedSystem_port_1_cast);

SharedReg299_out_to_MUX_Product226_impl_0_parent_implementedSystem_port_1_cast <= SharedReg299_out;
SharedReg331_out_to_MUX_Product226_impl_0_parent_implementedSystem_port_2_cast <= SharedReg331_out;
   MUX_Product226_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg299_out_to_MUX_Product226_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg331_out_to_MUX_Product226_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product226_impl_0_out);

   Delay1No330_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product226_impl_0_out,
                 Y => Delay1No330_out);

SharedReg232_out_to_MUX_Product226_impl_1_parent_implementedSystem_port_1_cast <= SharedReg232_out;
SharedReg233_out_to_MUX_Product226_impl_1_parent_implementedSystem_port_2_cast <= SharedReg233_out;
   MUX_Product226_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg232_out_to_MUX_Product226_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg233_out_to_MUX_Product226_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product226_impl_1_out);

   Delay1No331_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product226_impl_1_out,
                 Y => Delay1No331_out);

Delay1No332_out_to_Product326_impl_parent_implementedSystem_port_0_cast <= Delay1No332_out;
Delay1No333_out_to_Product326_impl_parent_implementedSystem_port_1_cast <= Delay1No333_out;
   Product326_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product326_impl_out,
                 X => Delay1No332_out_to_Product326_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No333_out_to_Product326_impl_parent_implementedSystem_port_1_cast);

SharedReg233_out_to_MUX_Product326_impl_0_parent_implementedSystem_port_1_cast <= SharedReg233_out;
SharedReg234_out_to_MUX_Product326_impl_0_parent_implementedSystem_port_2_cast <= SharedReg234_out;
   MUX_Product326_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg233_out_to_MUX_Product326_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg234_out_to_MUX_Product326_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product326_impl_0_out);

   Delay1No332_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product326_impl_0_out,
                 Y => Delay1No332_out);

SharedReg299_out_to_MUX_Product326_impl_1_parent_implementedSystem_port_1_cast <= SharedReg299_out;
SharedReg331_out_to_MUX_Product326_impl_1_parent_implementedSystem_port_2_cast <= SharedReg331_out;
   MUX_Product326_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg299_out_to_MUX_Product326_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg331_out_to_MUX_Product326_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product326_impl_1_out);

   Delay1No333_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product326_impl_1_out,
                 Y => Delay1No333_out);

Delay1No334_out_to_Subtract27_impl_parent_implementedSystem_port_0_cast <= Delay1No334_out;
Delay1No335_out_to_Subtract27_impl_parent_implementedSystem_port_1_cast <= Delay1No335_out;
   Subtract27_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract27_impl_out,
                 X => Delay1No334_out_to_Subtract27_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No335_out_to_Subtract27_impl_parent_implementedSystem_port_1_cast);

SharedReg191_out_to_MUX_Subtract27_impl_0_parent_implementedSystem_port_1_cast <= SharedReg191_out;
SharedReg122_out_to_MUX_Subtract27_impl_0_parent_implementedSystem_port_2_cast <= SharedReg122_out;
   MUX_Subtract27_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg191_out_to_MUX_Subtract27_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg122_out_to_MUX_Subtract27_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract27_impl_0_out);

   Delay1No334_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract27_impl_0_out,
                 Y => Delay1No334_out);

SharedReg194_out_to_MUX_Subtract27_impl_1_parent_implementedSystem_port_1_cast <= SharedReg194_out;
SharedReg127_out_to_MUX_Subtract27_impl_1_parent_implementedSystem_port_2_cast <= SharedReg127_out;
   MUX_Subtract27_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg194_out_to_MUX_Subtract27_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg127_out_to_MUX_Subtract27_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract27_impl_1_out);

   Delay1No335_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract27_impl_1_out,
                 Y => Delay1No335_out);

Delay1No336_out_to_Add83_impl_parent_implementedSystem_port_0_cast <= Delay1No336_out;
Delay1No337_out_to_Add83_impl_parent_implementedSystem_port_1_cast <= Delay1No337_out;
   Add83_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add83_impl_out,
                 X => Delay1No336_out_to_Add83_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No337_out_to_Add83_impl_parent_implementedSystem_port_1_cast);

SharedReg198_out_to_MUX_Add83_impl_0_parent_implementedSystem_port_1_cast <= SharedReg198_out;
SharedReg198_out_to_MUX_Add83_impl_0_parent_implementedSystem_port_2_cast <= SharedReg198_out;
   MUX_Add83_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg198_out_to_MUX_Add83_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg198_out_to_MUX_Add83_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add83_impl_0_out);

   Delay1No336_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add83_impl_0_out,
                 Y => Delay1No336_out);

SharedReg199_out_to_MUX_Add83_impl_1_parent_implementedSystem_port_1_cast <= SharedReg199_out;
SharedReg199_out_to_MUX_Add83_impl_1_parent_implementedSystem_port_2_cast <= SharedReg199_out;
   MUX_Add83_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg199_out_to_MUX_Add83_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg199_out_to_MUX_Add83_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add83_impl_1_out);

   Delay1No337_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add83_impl_1_out,
                 Y => Delay1No337_out);

Delay1No338_out_to_Product70_impl_parent_implementedSystem_port_0_cast <= Delay1No338_out;
Delay1No339_out_to_Product70_impl_parent_implementedSystem_port_1_cast <= Delay1No339_out;
   Product70_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product70_impl_out,
                 X => Delay1No338_out_to_Product70_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No339_out_to_Product70_impl_parent_implementedSystem_port_1_cast);

SharedReg342_out_to_MUX_Product70_impl_0_parent_implementedSystem_port_1_cast <= SharedReg342_out;
SharedReg336_out_to_MUX_Product70_impl_0_parent_implementedSystem_port_2_cast <= SharedReg336_out;
   MUX_Product70_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg342_out_to_MUX_Product70_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg336_out_to_MUX_Product70_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product70_impl_0_out);

   Delay1No338_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product70_impl_0_out,
                 Y => Delay1No338_out);

SharedReg70_out_to_MUX_Product70_impl_1_parent_implementedSystem_port_1_cast <= SharedReg70_out;
SharedReg65_out_to_MUX_Product70_impl_1_parent_implementedSystem_port_2_cast <= SharedReg65_out;
   MUX_Product70_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg70_out_to_MUX_Product70_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg65_out_to_MUX_Product70_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product70_impl_1_out);

   Delay1No339_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product70_impl_1_out,
                 Y => Delay1No339_out);

Delay1No340_out_to_Product142_impl_parent_implementedSystem_port_0_cast <= Delay1No340_out;
Delay1No341_out_to_Product142_impl_parent_implementedSystem_port_1_cast <= Delay1No341_out;
   Product142_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product142_impl_out,
                 X => Delay1No340_out_to_Product142_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No341_out_to_Product142_impl_parent_implementedSystem_port_1_cast);

SharedReg342_out_to_MUX_Product142_impl_0_parent_implementedSystem_port_1_cast <= SharedReg342_out;
SharedReg336_out_to_MUX_Product142_impl_0_parent_implementedSystem_port_2_cast <= SharedReg336_out;
   MUX_Product142_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg342_out_to_MUX_Product142_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg336_out_to_MUX_Product142_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product142_impl_0_out);

   Delay1No340_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product142_impl_0_out,
                 Y => Delay1No340_out);

SharedReg71_out_to_MUX_Product142_impl_1_parent_implementedSystem_port_1_cast <= SharedReg71_out;
SharedReg67_out_to_MUX_Product142_impl_1_parent_implementedSystem_port_2_cast <= SharedReg67_out;
   MUX_Product142_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg71_out_to_MUX_Product142_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg67_out_to_MUX_Product142_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product142_impl_1_out);

   Delay1No341_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product142_impl_1_out,
                 Y => Delay1No341_out);

Delay1No342_out_to_Product241_impl_parent_implementedSystem_port_0_cast <= Delay1No342_out;
Delay1No343_out_to_Product241_impl_parent_implementedSystem_port_1_cast <= Delay1No343_out;
   Product241_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product241_impl_out,
                 X => Delay1No342_out_to_Product241_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No343_out_to_Product241_impl_parent_implementedSystem_port_1_cast);

SharedReg343_out_to_MUX_Product241_impl_0_parent_implementedSystem_port_1_cast <= SharedReg343_out;
SharedReg337_out_to_MUX_Product241_impl_0_parent_implementedSystem_port_2_cast <= SharedReg337_out;
   MUX_Product241_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg343_out_to_MUX_Product241_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg337_out_to_MUX_Product241_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product241_impl_0_out);

   Delay1No342_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product241_impl_0_out,
                 Y => Delay1No342_out);

SharedReg70_out_to_MUX_Product241_impl_1_parent_implementedSystem_port_1_cast <= SharedReg70_out;
SharedReg65_out_to_MUX_Product241_impl_1_parent_implementedSystem_port_2_cast <= SharedReg65_out;
   MUX_Product241_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg70_out_to_MUX_Product241_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg65_out_to_MUX_Product241_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product241_impl_1_out);

   Delay1No343_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product241_impl_1_out,
                 Y => Delay1No343_out);

Delay1No344_out_to_Product341_impl_parent_implementedSystem_port_0_cast <= Delay1No344_out;
Delay1No345_out_to_Product341_impl_parent_implementedSystem_port_1_cast <= Delay1No345_out;
   Product341_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product341_impl_out,
                 X => Delay1No344_out_to_Product341_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No345_out_to_Product341_impl_parent_implementedSystem_port_1_cast);

SharedReg71_out_to_MUX_Product341_impl_0_parent_implementedSystem_port_1_cast <= SharedReg71_out;
SharedReg67_out_to_MUX_Product341_impl_0_parent_implementedSystem_port_2_cast <= SharedReg67_out;
   MUX_Product341_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg71_out_to_MUX_Product341_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg67_out_to_MUX_Product341_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product341_impl_0_out);

   Delay1No344_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product341_impl_0_out,
                 Y => Delay1No344_out);

SharedReg343_out_to_MUX_Product341_impl_1_parent_implementedSystem_port_1_cast <= SharedReg343_out;
SharedReg337_out_to_MUX_Product341_impl_1_parent_implementedSystem_port_2_cast <= SharedReg337_out;
   MUX_Product341_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg343_out_to_MUX_Product341_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg337_out_to_MUX_Product341_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product341_impl_1_out);

   Delay1No345_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product341_impl_1_out,
                 Y => Delay1No345_out);

Delay1No346_out_to_Subtract42_impl_parent_implementedSystem_port_0_cast <= Delay1No346_out;
Delay1No347_out_to_Subtract42_impl_parent_implementedSystem_port_1_cast <= Delay1No347_out;
   Subtract42_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract42_impl_out,
                 X => Delay1No346_out_to_Subtract42_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No347_out_to_Subtract42_impl_parent_implementedSystem_port_1_cast);

SharedReg166_out_to_MUX_Subtract42_impl_0_parent_implementedSystem_port_1_cast <= SharedReg166_out;
SharedReg197_out_to_MUX_Subtract42_impl_0_parent_implementedSystem_port_2_cast <= SharedReg197_out;
   MUX_Subtract42_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg166_out_to_MUX_Subtract42_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg197_out_to_MUX_Subtract42_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract42_impl_0_out);

   Delay1No346_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract42_impl_0_out,
                 Y => Delay1No346_out);

SharedReg172_out_to_MUX_Subtract42_impl_1_parent_implementedSystem_port_1_cast <= SharedReg172_out;
SharedReg200_out_to_MUX_Subtract42_impl_1_parent_implementedSystem_port_2_cast <= SharedReg200_out;
   MUX_Subtract42_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg172_out_to_MUX_Subtract42_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg200_out_to_MUX_Subtract42_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract42_impl_1_out);

   Delay1No347_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract42_impl_1_out,
                 Y => Delay1No347_out);

Delay1No348_out_to_Add84_impl_parent_implementedSystem_port_0_cast <= Delay1No348_out;
Delay1No349_out_to_Add84_impl_parent_implementedSystem_port_1_cast <= Delay1No349_out;
   Add84_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add84_impl_out,
                 X => Delay1No348_out_to_Add84_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No349_out_to_Add84_impl_parent_implementedSystem_port_1_cast);

SharedReg204_out_to_MUX_Add84_impl_0_parent_implementedSystem_port_1_cast <= SharedReg204_out;
SharedReg204_out_to_MUX_Add84_impl_0_parent_implementedSystem_port_2_cast <= SharedReg204_out;
   MUX_Add84_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg204_out_to_MUX_Add84_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg204_out_to_MUX_Add84_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add84_impl_0_out);

   Delay1No348_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add84_impl_0_out,
                 Y => Delay1No348_out);

SharedReg205_out_to_MUX_Add84_impl_1_parent_implementedSystem_port_1_cast <= SharedReg205_out;
SharedReg205_out_to_MUX_Add84_impl_1_parent_implementedSystem_port_2_cast <= SharedReg205_out;
   MUX_Add84_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg205_out_to_MUX_Add84_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg205_out_to_MUX_Add84_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add84_impl_1_out);

   Delay1No349_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add84_impl_1_out,
                 Y => Delay1No349_out);

Delay1No350_out_to_Product71_impl_parent_implementedSystem_port_0_cast <= Delay1No350_out;
Delay1No351_out_to_Product71_impl_parent_implementedSystem_port_1_cast <= Delay1No351_out;
   Product71_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product71_impl_out,
                 X => Delay1No350_out_to_Product71_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No351_out_to_Product71_impl_parent_implementedSystem_port_1_cast);

SharedReg346_out_to_MUX_Product71_impl_0_parent_implementedSystem_port_1_cast <= SharedReg346_out;
SharedReg340_out_to_MUX_Product71_impl_0_parent_implementedSystem_port_2_cast <= SharedReg340_out;
   MUX_Product71_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg346_out_to_MUX_Product71_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg340_out_to_MUX_Product71_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product71_impl_0_out);

   Delay1No350_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product71_impl_0_out,
                 Y => Delay1No350_out);

SharedReg72_out_to_MUX_Product71_impl_1_parent_implementedSystem_port_1_cast <= SharedReg72_out;
SharedReg236_out_to_MUX_Product71_impl_1_parent_implementedSystem_port_2_cast <= SharedReg236_out;
   MUX_Product71_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg72_out_to_MUX_Product71_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg236_out_to_MUX_Product71_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product71_impl_1_out);

   Delay1No351_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product71_impl_1_out,
                 Y => Delay1No351_out);

Delay1No352_out_to_Product143_impl_parent_implementedSystem_port_0_cast <= Delay1No352_out;
Delay1No353_out_to_Product143_impl_parent_implementedSystem_port_1_cast <= Delay1No353_out;
   Product143_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product143_impl_out,
                 X => Delay1No352_out_to_Product143_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No353_out_to_Product143_impl_parent_implementedSystem_port_1_cast);

SharedReg346_out_to_MUX_Product143_impl_0_parent_implementedSystem_port_1_cast <= SharedReg346_out;
SharedReg340_out_to_MUX_Product143_impl_0_parent_implementedSystem_port_2_cast <= SharedReg340_out;
   MUX_Product143_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg346_out_to_MUX_Product143_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg340_out_to_MUX_Product143_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product143_impl_0_out);

   Delay1No352_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product143_impl_0_out,
                 Y => Delay1No352_out);

SharedReg73_out_to_MUX_Product143_impl_1_parent_implementedSystem_port_1_cast <= SharedReg73_out;
SharedReg238_out_to_MUX_Product143_impl_1_parent_implementedSystem_port_2_cast <= SharedReg238_out;
   MUX_Product143_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg73_out_to_MUX_Product143_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg238_out_to_MUX_Product143_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product143_impl_1_out);

   Delay1No353_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product143_impl_1_out,
                 Y => Delay1No353_out);

Delay1No354_out_to_Product242_impl_parent_implementedSystem_port_0_cast <= Delay1No354_out;
Delay1No355_out_to_Product242_impl_parent_implementedSystem_port_1_cast <= Delay1No355_out;
   Product242_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product242_impl_out,
                 X => Delay1No354_out_to_Product242_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No355_out_to_Product242_impl_parent_implementedSystem_port_1_cast);

SharedReg347_out_to_MUX_Product242_impl_0_parent_implementedSystem_port_1_cast <= SharedReg347_out;
SharedReg341_out_to_MUX_Product242_impl_0_parent_implementedSystem_port_2_cast <= SharedReg341_out;
   MUX_Product242_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg347_out_to_MUX_Product242_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg341_out_to_MUX_Product242_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product242_impl_0_out);

   Delay1No354_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product242_impl_0_out,
                 Y => Delay1No354_out);

SharedReg72_out_to_MUX_Product242_impl_1_parent_implementedSystem_port_1_cast <= SharedReg72_out;
SharedReg236_out_to_MUX_Product242_impl_1_parent_implementedSystem_port_2_cast <= SharedReg236_out;
   MUX_Product242_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg72_out_to_MUX_Product242_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg236_out_to_MUX_Product242_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product242_impl_1_out);

   Delay1No355_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product242_impl_1_out,
                 Y => Delay1No355_out);

Delay1No356_out_to_Product342_impl_parent_implementedSystem_port_0_cast <= Delay1No356_out;
Delay1No357_out_to_Product342_impl_parent_implementedSystem_port_1_cast <= Delay1No357_out;
   Product342_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product342_impl_out,
                 X => Delay1No356_out_to_Product342_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No357_out_to_Product342_impl_parent_implementedSystem_port_1_cast);

SharedReg73_out_to_MUX_Product342_impl_0_parent_implementedSystem_port_1_cast <= SharedReg73_out;
SharedReg238_out_to_MUX_Product342_impl_0_parent_implementedSystem_port_2_cast <= SharedReg238_out;
   MUX_Product342_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg73_out_to_MUX_Product342_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg238_out_to_MUX_Product342_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product342_impl_0_out);

   Delay1No356_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product342_impl_0_out,
                 Y => Delay1No356_out);

SharedReg347_out_to_MUX_Product342_impl_1_parent_implementedSystem_port_1_cast <= SharedReg347_out;
SharedReg341_out_to_MUX_Product342_impl_1_parent_implementedSystem_port_2_cast <= SharedReg341_out;
   MUX_Product342_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg347_out_to_MUX_Product342_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg341_out_to_MUX_Product342_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product342_impl_1_out);

   Delay1No357_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product342_impl_1_out,
                 Y => Delay1No357_out);

Delay1No358_out_to_Subtract43_impl_parent_implementedSystem_port_0_cast <= Delay1No358_out;
Delay1No359_out_to_Subtract43_impl_parent_implementedSystem_port_1_cast <= Delay1No359_out;
   Subtract43_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract43_impl_out,
                 X => Delay1No358_out_to_Subtract43_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No359_out_to_Subtract43_impl_parent_implementedSystem_port_1_cast);

SharedReg129_out_to_MUX_Subtract43_impl_0_parent_implementedSystem_port_1_cast <= SharedReg129_out;
SharedReg203_out_to_MUX_Subtract43_impl_0_parent_implementedSystem_port_2_cast <= SharedReg203_out;
   MUX_Subtract43_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg129_out_to_MUX_Subtract43_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg203_out_to_MUX_Subtract43_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract43_impl_0_out);

   Delay1No358_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract43_impl_0_out,
                 Y => Delay1No358_out);

SharedReg135_out_to_MUX_Subtract43_impl_1_parent_implementedSystem_port_1_cast <= SharedReg135_out;
SharedReg206_out_to_MUX_Subtract43_impl_1_parent_implementedSystem_port_2_cast <= SharedReg206_out;
   MUX_Subtract43_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg135_out_to_MUX_Subtract43_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg206_out_to_MUX_Subtract43_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract43_impl_1_out);

   Delay1No359_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract43_impl_1_out,
                 Y => Delay1No359_out);

Delay1No360_out_to_Add85_impl_parent_implementedSystem_port_0_cast <= Delay1No360_out;
Delay1No361_out_to_Add85_impl_parent_implementedSystem_port_1_cast <= Delay1No361_out;
   Add85_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add85_impl_out,
                 X => Delay1No360_out_to_Add85_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No361_out_to_Add85_impl_parent_implementedSystem_port_1_cast);

SharedReg210_out_to_MUX_Add85_impl_0_parent_implementedSystem_port_1_cast <= SharedReg210_out;
SharedReg210_out_to_MUX_Add85_impl_0_parent_implementedSystem_port_2_cast <= SharedReg210_out;
   MUX_Add85_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg210_out_to_MUX_Add85_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg210_out_to_MUX_Add85_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add85_impl_0_out);

   Delay1No360_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add85_impl_0_out,
                 Y => Delay1No360_out);

SharedReg211_out_to_MUX_Add85_impl_1_parent_implementedSystem_port_1_cast <= SharedReg211_out;
SharedReg211_out_to_MUX_Add85_impl_1_parent_implementedSystem_port_2_cast <= SharedReg211_out;
   MUX_Add85_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg211_out_to_MUX_Add85_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg211_out_to_MUX_Add85_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add85_impl_1_out);

   Delay1No361_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add85_impl_1_out,
                 Y => Delay1No361_out);

Delay1No362_out_to_Product72_impl_parent_implementedSystem_port_0_cast <= Delay1No362_out;
Delay1No363_out_to_Product72_impl_parent_implementedSystem_port_1_cast <= Delay1No363_out;
   Product72_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product72_impl_out,
                 X => Delay1No362_out_to_Product72_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No363_out_to_Product72_impl_parent_implementedSystem_port_1_cast);

SharedReg348_out_to_MUX_Product72_impl_0_parent_implementedSystem_port_1_cast <= SharedReg348_out;
SharedReg338_out_to_MUX_Product72_impl_0_parent_implementedSystem_port_2_cast <= SharedReg338_out;
   MUX_Product72_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg348_out_to_MUX_Product72_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg338_out_to_MUX_Product72_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product72_impl_0_out);

   Delay1No362_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product72_impl_0_out,
                 Y => Delay1No362_out);

SharedReg224_out_to_MUX_Product72_impl_1_parent_implementedSystem_port_1_cast <= SharedReg224_out;
SharedReg239_out_to_MUX_Product72_impl_1_parent_implementedSystem_port_2_cast <= SharedReg239_out;
   MUX_Product72_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg224_out_to_MUX_Product72_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg239_out_to_MUX_Product72_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product72_impl_1_out);

   Delay1No363_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product72_impl_1_out,
                 Y => Delay1No363_out);

Delay1No364_out_to_Product144_impl_parent_implementedSystem_port_0_cast <= Delay1No364_out;
Delay1No365_out_to_Product144_impl_parent_implementedSystem_port_1_cast <= Delay1No365_out;
   Product144_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product144_impl_out,
                 X => Delay1No364_out_to_Product144_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No365_out_to_Product144_impl_parent_implementedSystem_port_1_cast);

SharedReg348_out_to_MUX_Product144_impl_0_parent_implementedSystem_port_1_cast <= SharedReg348_out;
SharedReg338_out_to_MUX_Product144_impl_0_parent_implementedSystem_port_2_cast <= SharedReg338_out;
   MUX_Product144_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg348_out_to_MUX_Product144_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg338_out_to_MUX_Product144_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product144_impl_0_out);

   Delay1No364_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product144_impl_0_out,
                 Y => Delay1No364_out);

SharedReg214_out_to_MUX_Product144_impl_1_parent_implementedSystem_port_1_cast <= SharedReg214_out;
SharedReg240_out_to_MUX_Product144_impl_1_parent_implementedSystem_port_2_cast <= SharedReg240_out;
   MUX_Product144_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg214_out_to_MUX_Product144_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg240_out_to_MUX_Product144_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product144_impl_1_out);

   Delay1No365_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product144_impl_1_out,
                 Y => Delay1No365_out);

Delay1No366_out_to_Product243_impl_parent_implementedSystem_port_0_cast <= Delay1No366_out;
Delay1No367_out_to_Product243_impl_parent_implementedSystem_port_1_cast <= Delay1No367_out;
   Product243_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product243_impl_out,
                 X => Delay1No366_out_to_Product243_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No367_out_to_Product243_impl_parent_implementedSystem_port_1_cast);

SharedReg349_out_to_MUX_Product243_impl_0_parent_implementedSystem_port_1_cast <= SharedReg349_out;
SharedReg339_out_to_MUX_Product243_impl_0_parent_implementedSystem_port_2_cast <= SharedReg339_out;
   MUX_Product243_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg349_out_to_MUX_Product243_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg339_out_to_MUX_Product243_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product243_impl_0_out);

   Delay1No366_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product243_impl_0_out,
                 Y => Delay1No366_out);

SharedReg224_out_to_MUX_Product243_impl_1_parent_implementedSystem_port_1_cast <= SharedReg224_out;
SharedReg239_out_to_MUX_Product243_impl_1_parent_implementedSystem_port_2_cast <= SharedReg239_out;
   MUX_Product243_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg224_out_to_MUX_Product243_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg239_out_to_MUX_Product243_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product243_impl_1_out);

   Delay1No367_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product243_impl_1_out,
                 Y => Delay1No367_out);

Delay1No368_out_to_Product343_impl_parent_implementedSystem_port_0_cast <= Delay1No368_out;
Delay1No369_out_to_Product343_impl_parent_implementedSystem_port_1_cast <= Delay1No369_out;
   Product343_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product343_impl_out,
                 X => Delay1No368_out_to_Product343_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No369_out_to_Product343_impl_parent_implementedSystem_port_1_cast);

SharedReg214_out_to_MUX_Product343_impl_0_parent_implementedSystem_port_1_cast <= SharedReg214_out;
SharedReg240_out_to_MUX_Product343_impl_0_parent_implementedSystem_port_2_cast <= SharedReg240_out;
   MUX_Product343_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg214_out_to_MUX_Product343_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg240_out_to_MUX_Product343_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product343_impl_0_out);

   Delay1No368_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product343_impl_0_out,
                 Y => Delay1No368_out);

SharedReg349_out_to_MUX_Product343_impl_1_parent_implementedSystem_port_1_cast <= SharedReg349_out;
SharedReg339_out_to_MUX_Product343_impl_1_parent_implementedSystem_port_2_cast <= SharedReg339_out;
   MUX_Product343_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg349_out_to_MUX_Product343_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg339_out_to_MUX_Product343_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product343_impl_1_out);

   Delay1No369_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product343_impl_1_out,
                 Y => Delay1No369_out);

Delay1No370_out_to_Subtract44_impl_parent_implementedSystem_port_0_cast <= Delay1No370_out;
Delay1No371_out_to_Subtract44_impl_parent_implementedSystem_port_1_cast <= Delay1No371_out;
   Subtract44_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract44_impl_out,
                 X => Delay1No370_out_to_Subtract44_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No371_out_to_Subtract44_impl_parent_implementedSystem_port_1_cast);

SharedReg118_out_to_MUX_Subtract44_impl_0_parent_implementedSystem_port_1_cast <= SharedReg118_out;
SharedReg209_out_to_MUX_Subtract44_impl_0_parent_implementedSystem_port_2_cast <= SharedReg209_out;
   MUX_Subtract44_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg118_out_to_MUX_Subtract44_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg209_out_to_MUX_Subtract44_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract44_impl_0_out);

   Delay1No370_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract44_impl_0_out,
                 Y => Delay1No370_out);

SharedReg130_out_to_MUX_Subtract44_impl_1_parent_implementedSystem_port_1_cast <= SharedReg130_out;
SharedReg212_out_to_MUX_Subtract44_impl_1_parent_implementedSystem_port_2_cast <= SharedReg212_out;
   MUX_Subtract44_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg130_out_to_MUX_Subtract44_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg212_out_to_MUX_Subtract44_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract44_impl_1_out);

   Delay1No371_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract44_impl_1_out,
                 Y => Delay1No371_out);

Delay1No372_out_to_Subtract45_impl_parent_implementedSystem_port_0_cast <= Delay1No372_out;
Delay1No373_out_to_Subtract45_impl_parent_implementedSystem_port_1_cast <= Delay1No373_out;
   Subtract45_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract45_impl_out,
                 X => Delay1No372_out_to_Subtract45_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No373_out_to_Subtract45_impl_parent_implementedSystem_port_1_cast);

SharedReg197_out_to_MUX_Subtract45_impl_0_parent_implementedSystem_port_1_cast <= SharedReg197_out;
SharedReg1_out_to_MUX_Subtract45_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1_out;
   MUX_Subtract45_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg197_out_to_MUX_Subtract45_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1_out_to_MUX_Subtract45_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract45_impl_0_out);

   Delay1No372_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract45_impl_0_out,
                 Y => Delay1No372_out);

SharedReg200_out_to_MUX_Subtract45_impl_1_parent_implementedSystem_port_1_cast <= SharedReg200_out;
SharedReg17_out_to_MUX_Subtract45_impl_1_parent_implementedSystem_port_2_cast <= SharedReg17_out;
   MUX_Subtract45_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg200_out_to_MUX_Subtract45_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg17_out_to_MUX_Subtract45_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract45_impl_1_out);

   Delay1No373_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract45_impl_1_out,
                 Y => Delay1No373_out);

Delay1No374_out_to_Add87_impl_parent_implementedSystem_port_0_cast <= Delay1No374_out;
Delay1No375_out_to_Add87_impl_parent_implementedSystem_port_1_cast <= Delay1No375_out;
   Add87_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add87_impl_out,
                 X => Delay1No374_out_to_Add87_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No375_out_to_Add87_impl_parent_implementedSystem_port_1_cast);

SharedReg217_out_to_MUX_Add87_impl_0_parent_implementedSystem_port_1_cast <= SharedReg217_out;
SharedReg217_out_to_MUX_Add87_impl_0_parent_implementedSystem_port_2_cast <= SharedReg217_out;
   MUX_Add87_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg217_out_to_MUX_Add87_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg217_out_to_MUX_Add87_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add87_impl_0_out);

   Delay1No374_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add87_impl_0_out,
                 Y => Delay1No374_out);

SharedReg218_out_to_MUX_Add87_impl_1_parent_implementedSystem_port_1_cast <= SharedReg218_out;
SharedReg218_out_to_MUX_Add87_impl_1_parent_implementedSystem_port_2_cast <= SharedReg218_out;
   MUX_Add87_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg218_out_to_MUX_Add87_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg218_out_to_MUX_Add87_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Add87_impl_1_out);

   Delay1No375_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add87_impl_1_out,
                 Y => Delay1No375_out);

Delay1No376_out_to_Product74_impl_parent_implementedSystem_port_0_cast <= Delay1No376_out;
Delay1No377_out_to_Product74_impl_parent_implementedSystem_port_1_cast <= Delay1No377_out;
   Product74_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product74_impl_out,
                 X => Delay1No376_out_to_Product74_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No377_out_to_Product74_impl_parent_implementedSystem_port_1_cast);

SharedReg350_out_to_MUX_Product74_impl_0_parent_implementedSystem_port_1_cast <= SharedReg350_out;
SharedReg344_out_to_MUX_Product74_impl_0_parent_implementedSystem_port_2_cast <= SharedReg344_out;
   MUX_Product74_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg350_out_to_MUX_Product74_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg344_out_to_MUX_Product74_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product74_impl_0_out);

   Delay1No376_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product74_impl_0_out,
                 Y => Delay1No376_out);

SharedReg221_out_to_MUX_Product74_impl_1_parent_implementedSystem_port_1_cast <= SharedReg221_out;
SharedReg64_out_to_MUX_Product74_impl_1_parent_implementedSystem_port_2_cast <= SharedReg64_out;
   MUX_Product74_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg221_out_to_MUX_Product74_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg64_out_to_MUX_Product74_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product74_impl_1_out);

   Delay1No377_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product74_impl_1_out,
                 Y => Delay1No377_out);

Delay1No378_out_to_Product146_impl_parent_implementedSystem_port_0_cast <= Delay1No378_out;
Delay1No379_out_to_Product146_impl_parent_implementedSystem_port_1_cast <= Delay1No379_out;
   Product146_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product146_impl_out,
                 X => Delay1No378_out_to_Product146_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No379_out_to_Product146_impl_parent_implementedSystem_port_1_cast);

SharedReg350_out_to_MUX_Product146_impl_0_parent_implementedSystem_port_1_cast <= SharedReg350_out;
SharedReg344_out_to_MUX_Product146_impl_0_parent_implementedSystem_port_2_cast <= SharedReg344_out;
   MUX_Product146_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg350_out_to_MUX_Product146_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg344_out_to_MUX_Product146_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product146_impl_0_out);

   Delay1No378_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product146_impl_0_out,
                 Y => Delay1No378_out);

SharedReg222_out_to_MUX_Product146_impl_1_parent_implementedSystem_port_1_cast <= SharedReg222_out;
SharedReg73_out_to_MUX_Product146_impl_1_parent_implementedSystem_port_2_cast <= SharedReg73_out;
   MUX_Product146_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg222_out_to_MUX_Product146_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg73_out_to_MUX_Product146_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product146_impl_1_out);

   Delay1No379_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product146_impl_1_out,
                 Y => Delay1No379_out);

Delay1No380_out_to_Product245_impl_parent_implementedSystem_port_0_cast <= Delay1No380_out;
Delay1No381_out_to_Product245_impl_parent_implementedSystem_port_1_cast <= Delay1No381_out;
   Product245_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product245_impl_out,
                 X => Delay1No380_out_to_Product245_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No381_out_to_Product245_impl_parent_implementedSystem_port_1_cast);

SharedReg351_out_to_MUX_Product245_impl_0_parent_implementedSystem_port_1_cast <= SharedReg351_out;
SharedReg345_out_to_MUX_Product245_impl_0_parent_implementedSystem_port_2_cast <= SharedReg345_out;
   MUX_Product245_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg351_out_to_MUX_Product245_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg345_out_to_MUX_Product245_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product245_impl_0_out);

   Delay1No380_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product245_impl_0_out,
                 Y => Delay1No380_out);

SharedReg221_out_to_MUX_Product245_impl_1_parent_implementedSystem_port_1_cast <= SharedReg221_out;
SharedReg64_out_to_MUX_Product245_impl_1_parent_implementedSystem_port_2_cast <= SharedReg64_out;
   MUX_Product245_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg221_out_to_MUX_Product245_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg64_out_to_MUX_Product245_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product245_impl_1_out);

   Delay1No381_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product245_impl_1_out,
                 Y => Delay1No381_out);

Delay1No382_out_to_Product345_impl_parent_implementedSystem_port_0_cast <= Delay1No382_out;
Delay1No383_out_to_Product345_impl_parent_implementedSystem_port_1_cast <= Delay1No383_out;
   Product345_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product345_impl_out,
                 X => Delay1No382_out_to_Product345_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No383_out_to_Product345_impl_parent_implementedSystem_port_1_cast);

SharedReg222_out_to_MUX_Product345_impl_0_parent_implementedSystem_port_1_cast <= SharedReg222_out;
SharedReg73_out_to_MUX_Product345_impl_0_parent_implementedSystem_port_2_cast <= SharedReg73_out;
   MUX_Product345_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg222_out_to_MUX_Product345_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg73_out_to_MUX_Product345_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product345_impl_0_out);

   Delay1No382_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product345_impl_0_out,
                 Y => Delay1No382_out);

SharedReg351_out_to_MUX_Product345_impl_1_parent_implementedSystem_port_1_cast <= SharedReg351_out;
SharedReg345_out_to_MUX_Product345_impl_1_parent_implementedSystem_port_2_cast <= SharedReg345_out;
   MUX_Product345_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg351_out_to_MUX_Product345_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg345_out_to_MUX_Product345_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Product345_impl_1_out);

   Delay1No383_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product345_impl_1_out,
                 Y => Delay1No383_out);

Delay1No384_out_to_Subtract46_impl_parent_implementedSystem_port_0_cast <= Delay1No384_out;
Delay1No385_out_to_Subtract46_impl_parent_implementedSystem_port_1_cast <= Delay1No385_out;
   Subtract46_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract46_impl_out,
                 X => Delay1No384_out_to_Subtract46_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No385_out_to_Subtract46_impl_parent_implementedSystem_port_1_cast);

SharedReg141_out_to_MUX_Subtract46_impl_0_parent_implementedSystem_port_1_cast <= SharedReg141_out;
SharedReg216_out_to_MUX_Subtract46_impl_0_parent_implementedSystem_port_2_cast <= SharedReg216_out;
   MUX_Subtract46_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg141_out_to_MUX_Subtract46_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg216_out_to_MUX_Subtract46_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract46_impl_0_out);

   Delay1No384_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract46_impl_0_out,
                 Y => Delay1No384_out);

SharedReg147_out_to_MUX_Subtract46_impl_1_parent_implementedSystem_port_1_cast <= SharedReg147_out;
SharedReg219_out_to_MUX_Subtract46_impl_1_parent_implementedSystem_port_2_cast <= SharedReg219_out;
   MUX_Subtract46_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg147_out_to_MUX_Subtract46_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg219_out_to_MUX_Subtract46_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract46_impl_1_out);

   Delay1No385_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract46_impl_1_out,
                 Y => Delay1No385_out);

Delay1No386_out_to_Subtract47_impl_parent_implementedSystem_port_0_cast <= Delay1No386_out;
Delay1No387_out_to_Subtract47_impl_parent_implementedSystem_port_1_cast <= Delay1No387_out;
   Subtract47_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract47_impl_out,
                 X => Delay1No386_out_to_Subtract47_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No387_out_to_Subtract47_impl_parent_implementedSystem_port_1_cast);

SharedReg203_out_to_MUX_Subtract47_impl_0_parent_implementedSystem_port_1_cast <= SharedReg203_out;
SharedReg2_out_to_MUX_Subtract47_impl_0_parent_implementedSystem_port_2_cast <= SharedReg2_out;
   MUX_Subtract47_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg203_out_to_MUX_Subtract47_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg2_out_to_MUX_Subtract47_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract47_impl_0_out);

   Delay1No386_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract47_impl_0_out,
                 Y => Delay1No386_out);

SharedReg206_out_to_MUX_Subtract47_impl_1_parent_implementedSystem_port_1_cast <= SharedReg206_out;
SharedReg18_out_to_MUX_Subtract47_impl_1_parent_implementedSystem_port_2_cast <= SharedReg18_out;
   MUX_Subtract47_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg206_out_to_MUX_Subtract47_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg18_out_to_MUX_Subtract47_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract47_impl_1_out);

   Delay1No387_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract47_impl_1_out,
                 Y => Delay1No387_out);

Delay1No388_out_to_Subtract48_impl_parent_implementedSystem_port_0_cast <= Delay1No388_out;
Delay1No389_out_to_Subtract48_impl_parent_implementedSystem_port_1_cast <= Delay1No389_out;
   Subtract48_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract48_impl_out,
                 X => Delay1No388_out_to_Subtract48_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No389_out_to_Subtract48_impl_parent_implementedSystem_port_1_cast);

SharedReg209_out_to_MUX_Subtract48_impl_0_parent_implementedSystem_port_1_cast <= SharedReg209_out;
SharedReg3_out_to_MUX_Subtract48_impl_0_parent_implementedSystem_port_2_cast <= SharedReg3_out;
   MUX_Subtract48_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg209_out_to_MUX_Subtract48_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg3_out_to_MUX_Subtract48_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract48_impl_0_out);

   Delay1No388_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract48_impl_0_out,
                 Y => Delay1No388_out);

SharedReg212_out_to_MUX_Subtract48_impl_1_parent_implementedSystem_port_1_cast <= SharedReg212_out;
SharedReg19_out_to_MUX_Subtract48_impl_1_parent_implementedSystem_port_2_cast <= SharedReg19_out;
   MUX_Subtract48_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg212_out_to_MUX_Subtract48_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg19_out_to_MUX_Subtract48_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract48_impl_1_out);

   Delay1No389_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract48_impl_1_out,
                 Y => Delay1No389_out);

Delay1No390_out_to_Subtract49_impl_parent_implementedSystem_port_0_cast <= Delay1No390_out;
Delay1No391_out_to_Subtract49_impl_parent_implementedSystem_port_1_cast <= Delay1No391_out;
   Subtract49_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract49_impl_out,
                 X => Delay1No390_out_to_Subtract49_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No391_out_to_Subtract49_impl_parent_implementedSystem_port_1_cast);

SharedReg216_out_to_MUX_Subtract49_impl_0_parent_implementedSystem_port_1_cast <= SharedReg216_out;
SharedReg183_out_to_MUX_Subtract49_impl_0_parent_implementedSystem_port_2_cast <= SharedReg183_out;
   MUX_Subtract49_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg216_out_to_MUX_Subtract49_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg183_out_to_MUX_Subtract49_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract49_impl_0_out);

   Delay1No390_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract49_impl_0_out,
                 Y => Delay1No390_out);

SharedReg219_out_to_MUX_Subtract49_impl_1_parent_implementedSystem_port_1_cast <= SharedReg219_out;
SharedReg221_out_to_MUX_Subtract49_impl_1_parent_implementedSystem_port_2_cast <= SharedReg221_out;
   MUX_Subtract49_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg219_out_to_MUX_Subtract49_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg221_out_to_MUX_Subtract49_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract49_impl_1_out);

   Delay1No391_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract49_impl_1_out,
                 Y => Delay1No391_out);

Delay1No392_out_to_Subtract50_impl_parent_implementedSystem_port_0_cast <= Delay1No392_out;
Delay1No393_out_to_Subtract50_impl_parent_implementedSystem_port_1_cast <= Delay1No393_out;
   Subtract50_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract50_impl_out,
                 X => Delay1No392_out_to_Subtract50_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No393_out_to_Subtract50_impl_parent_implementedSystem_port_1_cast);

SharedReg136_out_to_MUX_Subtract50_impl_0_parent_implementedSystem_port_1_cast <= SharedReg136_out;
SharedReg_out_to_MUX_Subtract50_impl_0_parent_implementedSystem_port_2_cast <= SharedReg_out;
   MUX_Subtract50_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg136_out_to_MUX_Subtract50_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg_out_to_MUX_Subtract50_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract50_impl_0_out);

   Delay1No392_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract50_impl_0_out,
                 Y => Delay1No392_out);

SharedReg142_out_to_MUX_Subtract50_impl_1_parent_implementedSystem_port_1_cast <= SharedReg142_out;
SharedReg16_out_to_MUX_Subtract50_impl_1_parent_implementedSystem_port_2_cast <= SharedReg16_out;
   MUX_Subtract50_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg142_out_to_MUX_Subtract50_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg16_out_to_MUX_Subtract50_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract50_impl_1_out);

   Delay1No393_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract50_impl_1_out,
                 Y => Delay1No393_out);

Delay1No394_out_to_Subtract52_impl_parent_implementedSystem_port_0_cast <= Delay1No394_out;
Delay1No395_out_to_Subtract52_impl_parent_implementedSystem_port_1_cast <= Delay1No395_out;
   Subtract52_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract52_impl_out,
                 X => Delay1No394_out_to_Subtract52_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No395_out_to_Subtract52_impl_parent_implementedSystem_port_1_cast);

SharedReg89_out_to_MUX_Subtract52_impl_0_parent_implementedSystem_port_1_cast <= SharedReg89_out;
SharedReg178_out_to_MUX_Subtract52_impl_0_parent_implementedSystem_port_2_cast <= SharedReg178_out;
   MUX_Subtract52_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg89_out_to_MUX_Subtract52_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg178_out_to_MUX_Subtract52_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract52_impl_0_out);

   Delay1No394_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract52_impl_0_out,
                 Y => Delay1No394_out);

SharedReg220_out_to_MUX_Subtract52_impl_1_parent_implementedSystem_port_1_cast <= SharedReg220_out;
SharedReg202_out_to_MUX_Subtract52_impl_1_parent_implementedSystem_port_2_cast <= SharedReg202_out;
   MUX_Subtract52_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg220_out_to_MUX_Subtract52_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg202_out_to_MUX_Subtract52_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract52_impl_1_out);

   Delay1No395_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract52_impl_1_out,
                 Y => Delay1No395_out);

Delay1No396_out_to_Subtract112_impl_parent_implementedSystem_port_0_cast <= Delay1No396_out;
Delay1No397_out_to_Subtract112_impl_parent_implementedSystem_port_1_cast <= Delay1No397_out;
   Subtract112_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract112_impl_out,
                 X => Delay1No396_out_to_Subtract112_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No397_out_to_Subtract112_impl_parent_implementedSystem_port_1_cast);

SharedReg90_out_to_MUX_Subtract112_impl_0_parent_implementedSystem_port_1_cast <= SharedReg90_out;
SharedReg222_out_to_MUX_Subtract112_impl_0_parent_implementedSystem_port_2_cast <= SharedReg222_out;
   MUX_Subtract112_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg90_out_to_MUX_Subtract112_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg222_out_to_MUX_Subtract112_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract112_impl_0_out);

   Delay1No396_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract112_impl_0_out,
                 Y => Delay1No396_out);

SharedReg215_out_to_MUX_Subtract112_impl_1_parent_implementedSystem_port_1_cast <= SharedReg215_out;
SharedReg99_out_to_MUX_Subtract112_impl_1_parent_implementedSystem_port_2_cast <= SharedReg99_out;
   MUX_Subtract112_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg215_out_to_MUX_Subtract112_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg99_out_to_MUX_Subtract112_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract112_impl_1_out);

   Delay1No397_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract112_impl_1_out,
                 Y => Delay1No397_out);

Delay1No398_out_to_Subtract114_impl_parent_implementedSystem_port_0_cast <= Delay1No398_out;
Delay1No399_out_to_Subtract114_impl_parent_implementedSystem_port_1_cast <= Delay1No399_out;
   Subtract114_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract114_impl_out,
                 X => Delay1No398_out_to_Subtract114_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No399_out_to_Subtract114_impl_parent_implementedSystem_port_1_cast);

SharedReg83_out_to_MUX_Subtract114_impl_0_parent_implementedSystem_port_1_cast <= SharedReg83_out;
SharedReg208_out_to_MUX_Subtract114_impl_0_parent_implementedSystem_port_2_cast <= SharedReg208_out;
   MUX_Subtract114_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg83_out_to_MUX_Subtract114_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg208_out_to_MUX_Subtract114_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract114_impl_0_out);

   Delay1No398_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract114_impl_0_out,
                 Y => Delay1No398_out);

SharedReg123_out_to_MUX_Subtract114_impl_1_parent_implementedSystem_port_1_cast <= SharedReg123_out;
SharedReg94_out_to_MUX_Subtract114_impl_1_parent_implementedSystem_port_2_cast <= SharedReg94_out;
   MUX_Subtract114_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg123_out_to_MUX_Subtract114_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg94_out_to_MUX_Subtract114_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract114_impl_1_out);

   Delay1No399_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract114_impl_1_out,
                 Y => Delay1No399_out);

Delay1No400_out_to_Subtract55_impl_parent_implementedSystem_port_0_cast <= Delay1No400_out;
Delay1No401_out_to_Subtract55_impl_parent_implementedSystem_port_1_cast <= Delay1No401_out;
   Subtract55_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract55_impl_out,
                 X => Delay1No400_out_to_Subtract55_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No401_out_to_Subtract55_impl_parent_implementedSystem_port_1_cast);

SharedReg84_out_to_MUX_Subtract55_impl_0_parent_implementedSystem_port_1_cast <= SharedReg84_out;
SharedReg223_out_to_MUX_Subtract55_impl_0_parent_implementedSystem_port_2_cast <= SharedReg223_out;
   MUX_Subtract55_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg84_out_to_MUX_Subtract55_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg223_out_to_MUX_Subtract55_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract55_impl_0_out);

   Delay1No400_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract55_impl_0_out,
                 Y => Delay1No400_out);

SharedReg124_out_to_MUX_Subtract55_impl_1_parent_implementedSystem_port_1_cast <= SharedReg124_out;
SharedReg105_out_to_MUX_Subtract55_impl_1_parent_implementedSystem_port_2_cast <= SharedReg105_out;
   MUX_Subtract55_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg124_out_to_MUX_Subtract55_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg105_out_to_MUX_Subtract55_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract55_impl_1_out);

   Delay1No401_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract55_impl_1_out,
                 Y => Delay1No401_out);

Delay1No402_out_to_Subtract115_impl_parent_implementedSystem_port_0_cast <= Delay1No402_out;
Delay1No403_out_to_Subtract115_impl_parent_implementedSystem_port_1_cast <= Delay1No403_out;
   Subtract115_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract115_impl_out,
                 X => Delay1No402_out_to_Subtract115_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No403_out_to_Subtract115_impl_parent_implementedSystem_port_1_cast);

SharedReg99_out_to_MUX_Subtract115_impl_0_parent_implementedSystem_port_1_cast <= SharedReg99_out;
SharedReg215_out_to_MUX_Subtract115_impl_0_parent_implementedSystem_port_2_cast <= SharedReg215_out;
   MUX_Subtract115_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg99_out_to_MUX_Subtract115_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg215_out_to_MUX_Subtract115_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract115_impl_0_out);

   Delay1No402_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract115_impl_0_out,
                 Y => Delay1No402_out);

SharedReg105_out_to_MUX_Subtract115_impl_1_parent_implementedSystem_port_1_cast <= SharedReg105_out;
SharedReg100_out_to_MUX_Subtract115_impl_1_parent_implementedSystem_port_2_cast <= SharedReg100_out;
   MUX_Subtract115_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg105_out_to_MUX_Subtract115_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg100_out_to_MUX_Subtract115_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract115_impl_1_out);

   Delay1No403_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract115_impl_1_out,
                 Y => Delay1No403_out);

Delay1No404_out_to_Subtract56_impl_parent_implementedSystem_port_0_cast <= Delay1No404_out;
Delay1No405_out_to_Subtract56_impl_parent_implementedSystem_port_1_cast <= Delay1No405_out;
   Subtract56_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract56_impl_out,
                 X => Delay1No404_out_to_Subtract56_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No405_out_to_Subtract56_impl_parent_implementedSystem_port_1_cast);

SharedReg94_out_to_MUX_Subtract56_impl_0_parent_implementedSystem_port_1_cast <= SharedReg94_out;
SharedReg89_out_to_MUX_Subtract56_impl_0_parent_implementedSystem_port_2_cast <= SharedReg89_out;
   MUX_Subtract56_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg94_out_to_MUX_Subtract56_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg89_out_to_MUX_Subtract56_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract56_impl_0_out);

   Delay1No404_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract56_impl_0_out,
                 Y => Delay1No404_out);

SharedReg100_out_to_MUX_Subtract56_impl_1_parent_implementedSystem_port_1_cast <= SharedReg100_out;
SharedReg111_out_to_MUX_Subtract56_impl_1_parent_implementedSystem_port_2_cast <= SharedReg111_out;
   MUX_Subtract56_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg100_out_to_MUX_Subtract56_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg111_out_to_MUX_Subtract56_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract56_impl_1_out);

   Delay1No405_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract56_impl_1_out,
                 Y => Delay1No405_out);

Delay1No406_out_to_Subtract116_impl_parent_implementedSystem_port_0_cast <= Delay1No406_out;
Delay1No407_out_to_Subtract116_impl_parent_implementedSystem_port_1_cast <= Delay1No407_out;
   Subtract116_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract116_impl_out,
                 X => Delay1No406_out_to_Subtract116_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No407_out_to_Subtract116_impl_parent_implementedSystem_port_1_cast);

Delay2No49_out_to_MUX_Subtract116_impl_0_parent_implementedSystem_port_1_cast <= Delay2No49_out;
SharedReg84_out_to_MUX_Subtract116_impl_0_parent_implementedSystem_port_2_cast <= SharedReg84_out;
   MUX_Subtract116_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No49_out_to_MUX_Subtract116_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg84_out_to_MUX_Subtract116_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract116_impl_0_out);

   Delay1No406_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract116_impl_0_out,
                 Y => Delay1No406_out);

Delay2No51_out_to_MUX_Subtract116_impl_1_parent_implementedSystem_port_1_cast <= Delay2No51_out;
SharedReg106_out_to_MUX_Subtract116_impl_1_parent_implementedSystem_port_2_cast <= SharedReg106_out;
   MUX_Subtract116_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No51_out_to_MUX_Subtract116_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg106_out_to_MUX_Subtract116_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract116_impl_1_out);

   Delay1No407_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract116_impl_1_out,
                 Y => Delay1No407_out);

Delay1No408_out_to_Subtract57_impl_parent_implementedSystem_port_0_cast <= Delay1No408_out;
Delay1No409_out_to_Subtract57_impl_parent_implementedSystem_port_1_cast <= Delay1No409_out;
   Subtract57_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract57_impl_out,
                 X => Delay1No408_out_to_Subtract57_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No409_out_to_Subtract57_impl_parent_implementedSystem_port_1_cast);

Delay2No48_out_to_MUX_Subtract57_impl_0_parent_implementedSystem_port_1_cast <= Delay2No48_out;
SharedReg81_out_to_MUX_Subtract57_impl_0_parent_implementedSystem_port_2_cast <= SharedReg81_out;
   MUX_Subtract57_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No48_out_to_MUX_Subtract57_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg81_out_to_MUX_Subtract57_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract57_impl_0_out);

   Delay1No408_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract57_impl_0_out,
                 Y => Delay1No408_out);

Delay2No50_out_to_MUX_Subtract57_impl_1_parent_implementedSystem_port_1_cast <= Delay2No50_out;
SharedReg117_out_to_MUX_Subtract57_impl_1_parent_implementedSystem_port_2_cast <= SharedReg117_out;
   MUX_Subtract57_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No50_out_to_MUX_Subtract57_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg117_out_to_MUX_Subtract57_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract57_impl_1_out);

   Delay1No409_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract57_impl_1_out,
                 Y => Delay1No409_out);

Delay1No410_out_to_Subtract117_impl_parent_implementedSystem_port_0_cast <= Delay1No410_out;
Delay1No411_out_to_Subtract117_impl_parent_implementedSystem_port_1_cast <= Delay1No411_out;
   Subtract117_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract117_impl_out,
                 X => Delay1No410_out_to_Subtract117_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No411_out_to_Subtract117_impl_parent_implementedSystem_port_1_cast);

Delay2No41_out_to_MUX_Subtract117_impl_0_parent_implementedSystem_port_1_cast <= Delay2No41_out;
SharedReg90_out_to_MUX_Subtract117_impl_0_parent_implementedSystem_port_2_cast <= SharedReg90_out;
   MUX_Subtract117_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No41_out_to_MUX_Subtract117_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg90_out_to_MUX_Subtract117_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract117_impl_0_out);

   Delay1No410_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract117_impl_0_out,
                 Y => Delay1No410_out);

Delay2No43_out_to_MUX_Subtract117_impl_1_parent_implementedSystem_port_1_cast <= Delay2No43_out;
SharedReg112_out_to_MUX_Subtract117_impl_1_parent_implementedSystem_port_2_cast <= SharedReg112_out;
   MUX_Subtract117_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No43_out_to_MUX_Subtract117_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg112_out_to_MUX_Subtract117_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract117_impl_1_out);

   Delay1No411_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract117_impl_1_out,
                 Y => Delay1No411_out);

Delay1No412_out_to_Subtract59_impl_parent_implementedSystem_port_0_cast <= Delay1No412_out;
Delay1No413_out_to_Subtract59_impl_parent_implementedSystem_port_1_cast <= Delay1No413_out;
   Subtract59_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract59_impl_out,
                 X => Delay1No412_out_to_Subtract59_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No413_out_to_Subtract59_impl_parent_implementedSystem_port_1_cast);

Delay2No40_out_to_MUX_Subtract59_impl_0_parent_implementedSystem_port_1_cast <= Delay2No40_out;
SharedReg123_out_to_MUX_Subtract59_impl_0_parent_implementedSystem_port_2_cast <= SharedReg123_out;
   MUX_Subtract59_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No40_out_to_MUX_Subtract59_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg123_out_to_MUX_Subtract59_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract59_impl_0_out);

   Delay1No412_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract59_impl_0_out,
                 Y => Delay1No412_out);

Delay2No42_out_to_MUX_Subtract59_impl_1_parent_implementedSystem_port_1_cast <= Delay2No42_out;
SharedReg165_out_to_MUX_Subtract59_impl_1_parent_implementedSystem_port_2_cast <= SharedReg165_out;
   MUX_Subtract59_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No42_out_to_MUX_Subtract59_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg165_out_to_MUX_Subtract59_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract59_impl_1_out);

   Delay1No413_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract59_impl_1_out,
                 Y => Delay1No413_out);

Delay1No414_out_to_Subtract119_impl_parent_implementedSystem_port_0_cast <= Delay1No414_out;
Delay1No415_out_to_Subtract119_impl_parent_implementedSystem_port_1_cast <= Delay1No415_out;
   Subtract119_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract119_impl_out,
                 X => Delay1No414_out_to_Subtract119_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No415_out_to_Subtract119_impl_parent_implementedSystem_port_1_cast);

Delay2No45_out_to_MUX_Subtract119_impl_0_parent_implementedSystem_port_1_cast <= Delay2No45_out;
SharedReg118_out_to_MUX_Subtract119_impl_0_parent_implementedSystem_port_2_cast <= SharedReg118_out;
   MUX_Subtract119_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No45_out_to_MUX_Subtract119_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg118_out_to_MUX_Subtract119_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract119_impl_0_out);

   Delay1No414_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract119_impl_0_out,
                 Y => Delay1No414_out);

Delay2No53_out_to_MUX_Subtract119_impl_1_parent_implementedSystem_port_1_cast <= Delay2No53_out;
SharedReg160_out_to_MUX_Subtract119_impl_1_parent_implementedSystem_port_2_cast <= SharedReg160_out;
   MUX_Subtract119_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No53_out_to_MUX_Subtract119_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg160_out_to_MUX_Subtract119_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract119_impl_1_out);

   Delay1No415_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract119_impl_1_out,
                 Y => Delay1No415_out);

Delay1No416_out_to_Subtract62_impl_parent_implementedSystem_port_0_cast <= Delay1No416_out;
Delay1No417_out_to_Subtract62_impl_parent_implementedSystem_port_1_cast <= Delay1No417_out;
   Subtract62_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract62_impl_out,
                 X => Delay1No416_out_to_Subtract62_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No417_out_to_Subtract62_impl_parent_implementedSystem_port_1_cast);

Delay2No44_out_to_MUX_Subtract62_impl_0_parent_implementedSystem_port_1_cast <= Delay2No44_out;
SharedReg4_out_to_MUX_Subtract62_impl_0_parent_implementedSystem_port_2_cast <= SharedReg4_out;
   MUX_Subtract62_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No44_out_to_MUX_Subtract62_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg4_out_to_MUX_Subtract62_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract62_impl_0_out);

   Delay1No416_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract62_impl_0_out,
                 Y => Delay1No416_out);

Delay2No52_out_to_MUX_Subtract62_impl_1_parent_implementedSystem_port_1_cast <= Delay2No52_out;
SharedReg20_out_to_MUX_Subtract62_impl_1_parent_implementedSystem_port_2_cast <= SharedReg20_out;
   MUX_Subtract62_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No52_out_to_MUX_Subtract62_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg20_out_to_MUX_Subtract62_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract62_impl_1_out);

   Delay1No417_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract62_impl_1_out,
                 Y => Delay1No417_out);

Delay1No418_out_to_Subtract122_impl_parent_implementedSystem_port_0_cast <= Delay1No418_out;
Delay1No419_out_to_Subtract122_impl_parent_implementedSystem_port_1_cast <= Delay1No419_out;
   Subtract122_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract122_impl_out,
                 X => Delay1No418_out_to_Subtract122_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No419_out_to_Subtract122_impl_parent_implementedSystem_port_1_cast);

Delay2No47_out_to_MUX_Subtract122_impl_0_parent_implementedSystem_port_1_cast <= Delay2No47_out;
SharedReg5_out_to_MUX_Subtract122_impl_0_parent_implementedSystem_port_2_cast <= SharedReg5_out;
   MUX_Subtract122_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No47_out_to_MUX_Subtract122_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg5_out_to_MUX_Subtract122_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract122_impl_0_out);

   Delay1No418_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract122_impl_0_out,
                 Y => Delay1No418_out);

Delay2No55_out_to_MUX_Subtract122_impl_1_parent_implementedSystem_port_1_cast <= Delay2No55_out;
SharedReg21_out_to_MUX_Subtract122_impl_1_parent_implementedSystem_port_2_cast <= SharedReg21_out;
   MUX_Subtract122_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No55_out_to_MUX_Subtract122_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg21_out_to_MUX_Subtract122_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract122_impl_1_out);

   Delay1No419_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract122_impl_1_out,
                 Y => Delay1No419_out);

Delay1No420_out_to_Subtract63_impl_parent_implementedSystem_port_0_cast <= Delay1No420_out;
Delay1No421_out_to_Subtract63_impl_parent_implementedSystem_port_1_cast <= Delay1No421_out;
   Subtract63_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract63_impl_out,
                 X => Delay1No420_out_to_Subtract63_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No421_out_to_Subtract63_impl_parent_implementedSystem_port_1_cast);

Delay2No46_out_to_MUX_Subtract63_impl_0_parent_implementedSystem_port_1_cast <= Delay2No46_out;
SharedReg129_out_to_MUX_Subtract63_impl_0_parent_implementedSystem_port_2_cast <= SharedReg129_out;
   MUX_Subtract63_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No46_out_to_MUX_Subtract63_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg129_out_to_MUX_Subtract63_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract63_impl_0_out);

   Delay1No420_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract63_impl_0_out,
                 Y => Delay1No420_out);

Delay2No54_out_to_MUX_Subtract63_impl_1_parent_implementedSystem_port_1_cast <= Delay2No54_out;
SharedReg141_out_to_MUX_Subtract63_impl_1_parent_implementedSystem_port_2_cast <= SharedReg141_out;
   MUX_Subtract63_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No54_out_to_MUX_Subtract63_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg141_out_to_MUX_Subtract63_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract63_impl_1_out);

   Delay1No421_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract63_impl_1_out,
                 Y => Delay1No421_out);

Delay1No422_out_to_Subtract123_impl_parent_implementedSystem_port_0_cast <= Delay1No422_out;
Delay1No423_out_to_Subtract123_impl_parent_implementedSystem_port_1_cast <= Delay1No423_out;
   Subtract123_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract123_impl_out,
                 X => Delay1No422_out_to_Subtract123_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No423_out_to_Subtract123_impl_parent_implementedSystem_port_1_cast);

SharedReg111_out_to_MUX_Subtract123_impl_0_parent_implementedSystem_port_1_cast <= SharedReg111_out;
SharedReg124_out_to_MUX_Subtract123_impl_0_parent_implementedSystem_port_2_cast <= SharedReg124_out;
   MUX_Subtract123_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg111_out_to_MUX_Subtract123_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg124_out_to_MUX_Subtract123_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract123_impl_0_out);

   Delay1No422_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract123_impl_0_out,
                 Y => Delay1No422_out);

SharedReg117_out_to_MUX_Subtract123_impl_1_parent_implementedSystem_port_1_cast <= SharedReg117_out;
SharedReg136_out_to_MUX_Subtract123_impl_1_parent_implementedSystem_port_2_cast <= SharedReg136_out;
   MUX_Subtract123_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg117_out_to_MUX_Subtract123_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg136_out_to_MUX_Subtract123_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract123_impl_1_out);

   Delay1No423_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract123_impl_1_out,
                 Y => Delay1No423_out);

Delay1No424_out_to_Subtract127_impl_parent_implementedSystem_port_0_cast <= Delay1No424_out;
Delay1No425_out_to_Subtract127_impl_parent_implementedSystem_port_1_cast <= Delay1No425_out;
   Subtract127_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract127_impl_out,
                 X => Delay1No424_out_to_Subtract127_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No425_out_to_Subtract127_impl_parent_implementedSystem_port_1_cast);

SharedReg106_out_to_MUX_Subtract127_impl_0_parent_implementedSystem_port_1_cast <= SharedReg106_out;
SharedReg6_out_to_MUX_Subtract127_impl_0_parent_implementedSystem_port_2_cast <= SharedReg6_out;
   MUX_Subtract127_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg106_out_to_MUX_Subtract127_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg6_out_to_MUX_Subtract127_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract127_impl_0_out);

   Delay1No424_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract127_impl_0_out,
                 Y => Delay1No424_out);

SharedReg112_out_to_MUX_Subtract127_impl_1_parent_implementedSystem_port_1_cast <= SharedReg112_out;
SharedReg22_out_to_MUX_Subtract127_impl_1_parent_implementedSystem_port_2_cast <= SharedReg22_out;
   MUX_Subtract127_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg112_out_to_MUX_Subtract127_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg22_out_to_MUX_Subtract127_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract127_impl_1_out);

   Delay1No425_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract127_impl_1_out,
                 Y => Delay1No425_out);

Delay1No426_out_to_Subtract68_impl_parent_implementedSystem_port_0_cast <= Delay1No426_out;
Delay1No427_out_to_Subtract68_impl_parent_implementedSystem_port_1_cast <= Delay1No427_out;
   Subtract68_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract68_impl_out,
                 X => Delay1No426_out_to_Subtract68_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No427_out_to_Subtract68_impl_parent_implementedSystem_port_1_cast);

SharedReg171_out_to_MUX_Subtract68_impl_0_parent_implementedSystem_port_1_cast <= SharedReg171_out;
SharedReg7_out_to_MUX_Subtract68_impl_0_parent_implementedSystem_port_2_cast <= SharedReg7_out;
   MUX_Subtract68_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg171_out_to_MUX_Subtract68_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg7_out_to_MUX_Subtract68_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract68_impl_0_out);

   Delay1No426_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract68_impl_0_out,
                 Y => Delay1No426_out);

SharedReg177_out_to_MUX_Subtract68_impl_1_parent_implementedSystem_port_1_cast <= SharedReg177_out;
SharedReg23_out_to_MUX_Subtract68_impl_1_parent_implementedSystem_port_2_cast <= SharedReg23_out;
   MUX_Subtract68_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg177_out_to_MUX_Subtract68_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg23_out_to_MUX_Subtract68_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract68_impl_1_out);

   Delay1No427_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract68_impl_1_out,
                 Y => Delay1No427_out);

Delay1No428_out_to_Subtract71_impl_parent_implementedSystem_port_0_cast <= Delay1No428_out;
Delay1No429_out_to_Subtract71_impl_parent_implementedSystem_port_1_cast <= Delay1No429_out;
   Subtract71_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract71_impl_out,
                 X => Delay1No428_out_to_Subtract71_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No429_out_to_Subtract71_impl_parent_implementedSystem_port_1_cast);

SharedReg153_out_to_MUX_Subtract71_impl_0_parent_implementedSystem_port_1_cast <= SharedReg153_out;
SharedReg8_out_to_MUX_Subtract71_impl_0_parent_implementedSystem_port_2_cast <= SharedReg8_out;
   MUX_Subtract71_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg153_out_to_MUX_Subtract71_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg8_out_to_MUX_Subtract71_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract71_impl_0_out);

   Delay1No428_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract71_impl_0_out,
                 Y => Delay1No428_out);

SharedReg159_out_to_MUX_Subtract71_impl_1_parent_implementedSystem_port_1_cast <= SharedReg159_out;
SharedReg24_out_to_MUX_Subtract71_impl_1_parent_implementedSystem_port_2_cast <= SharedReg24_out;
   MUX_Subtract71_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg159_out_to_MUX_Subtract71_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg24_out_to_MUX_Subtract71_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract71_impl_1_out);

   Delay1No429_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract71_impl_1_out,
                 Y => Delay1No429_out);

Delay1No430_out_to_Subtract131_impl_parent_implementedSystem_port_0_cast <= Delay1No430_out;
Delay1No431_out_to_Subtract131_impl_parent_implementedSystem_port_1_cast <= Delay1No431_out;
   Subtract131_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract131_impl_out,
                 X => Delay1No430_out_to_Subtract131_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No431_out_to_Subtract131_impl_parent_implementedSystem_port_1_cast);

SharedReg148_out_to_MUX_Subtract131_impl_0_parent_implementedSystem_port_1_cast <= SharedReg148_out;
SharedReg9_out_to_MUX_Subtract131_impl_0_parent_implementedSystem_port_2_cast <= SharedReg9_out;
   MUX_Subtract131_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg148_out_to_MUX_Subtract131_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg9_out_to_MUX_Subtract131_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract131_impl_0_out);

   Delay1No430_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract131_impl_0_out,
                 Y => Delay1No430_out);

SharedReg154_out_to_MUX_Subtract131_impl_1_parent_implementedSystem_port_1_cast <= SharedReg154_out;
SharedReg25_out_to_MUX_Subtract131_impl_1_parent_implementedSystem_port_2_cast <= SharedReg25_out;
   MUX_Subtract131_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg154_out_to_MUX_Subtract131_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg25_out_to_MUX_Subtract131_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract131_impl_1_out);

   Delay1No431_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract131_impl_1_out,
                 Y => Delay1No431_out);

Delay1No432_out_to_Subtract72_impl_parent_implementedSystem_port_0_cast <= Delay1No432_out;
Delay1No433_out_to_Subtract72_impl_parent_implementedSystem_port_1_cast <= Delay1No433_out;
   Subtract72_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract72_impl_out,
                 X => Delay1No432_out_to_Subtract72_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No433_out_to_Subtract72_impl_parent_implementedSystem_port_1_cast);

SharedReg183_out_to_MUX_Subtract72_impl_0_parent_implementedSystem_port_1_cast <= SharedReg183_out;
SharedReg10_out_to_MUX_Subtract72_impl_0_parent_implementedSystem_port_2_cast <= SharedReg10_out;
   MUX_Subtract72_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg183_out_to_MUX_Subtract72_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg10_out_to_MUX_Subtract72_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract72_impl_0_out);

   Delay1No432_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract72_impl_0_out,
                 Y => Delay1No432_out);

SharedReg189_out_to_MUX_Subtract72_impl_1_parent_implementedSystem_port_1_cast <= SharedReg189_out;
SharedReg26_out_to_MUX_Subtract72_impl_1_parent_implementedSystem_port_2_cast <= SharedReg26_out;
   MUX_Subtract72_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg189_out_to_MUX_Subtract72_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg26_out_to_MUX_Subtract72_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract72_impl_1_out);

   Delay1No433_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract72_impl_1_out,
                 Y => Delay1No433_out);

Delay1No434_out_to_Subtract132_impl_parent_implementedSystem_port_0_cast <= Delay1No434_out;
Delay1No435_out_to_Subtract132_impl_parent_implementedSystem_port_1_cast <= Delay1No435_out;
   Subtract132_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract132_impl_out,
                 X => Delay1No434_out_to_Subtract132_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No435_out_to_Subtract132_impl_parent_implementedSystem_port_1_cast);

SharedReg178_out_to_MUX_Subtract132_impl_0_parent_implementedSystem_port_1_cast <= SharedReg178_out;
SharedReg11_out_to_MUX_Subtract132_impl_0_parent_implementedSystem_port_2_cast <= SharedReg11_out;
   MUX_Subtract132_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg178_out_to_MUX_Subtract132_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg11_out_to_MUX_Subtract132_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract132_impl_0_out);

   Delay1No434_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract132_impl_0_out,
                 Y => Delay1No434_out);

SharedReg184_out_to_MUX_Subtract132_impl_1_parent_implementedSystem_port_1_cast <= SharedReg184_out;
SharedReg27_out_to_MUX_Subtract132_impl_1_parent_implementedSystem_port_2_cast <= SharedReg27_out;
   MUX_Subtract132_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg184_out_to_MUX_Subtract132_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg27_out_to_MUX_Subtract132_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract132_impl_1_out);

   Delay1No435_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract132_impl_1_out,
                 Y => Delay1No435_out);

Delay1No436_out_to_Subtract74_impl_parent_implementedSystem_port_0_cast <= Delay1No436_out;
Delay1No437_out_to_Subtract74_impl_parent_implementedSystem_port_1_cast <= Delay1No437_out;
   Subtract74_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract74_impl_out,
                 X => Delay1No436_out_to_Subtract74_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No437_out_to_Subtract74_impl_parent_implementedSystem_port_1_cast);

SharedReg195_out_to_MUX_Subtract74_impl_0_parent_implementedSystem_port_1_cast <= SharedReg195_out;
SharedReg12_out_to_MUX_Subtract74_impl_0_parent_implementedSystem_port_2_cast <= SharedReg12_out;
   MUX_Subtract74_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg195_out_to_MUX_Subtract74_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg12_out_to_MUX_Subtract74_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract74_impl_0_out);

   Delay1No436_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract74_impl_0_out,
                 Y => Delay1No436_out);

SharedReg201_out_to_MUX_Subtract74_impl_1_parent_implementedSystem_port_1_cast <= SharedReg201_out;
SharedReg28_out_to_MUX_Subtract74_impl_1_parent_implementedSystem_port_2_cast <= SharedReg28_out;
   MUX_Subtract74_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg201_out_to_MUX_Subtract74_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg28_out_to_MUX_Subtract74_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract74_impl_1_out);

   Delay1No437_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract74_impl_1_out,
                 Y => Delay1No437_out);

Delay1No438_out_to_Subtract134_impl_parent_implementedSystem_port_0_cast <= Delay1No438_out;
Delay1No439_out_to_Subtract134_impl_parent_implementedSystem_port_1_cast <= Delay1No439_out;
   Subtract134_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract134_impl_out,
                 X => Delay1No438_out_to_Subtract134_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No439_out_to_Subtract134_impl_parent_implementedSystem_port_1_cast);

SharedReg190_out_to_MUX_Subtract134_impl_0_parent_implementedSystem_port_1_cast <= SharedReg190_out;
SharedReg13_out_to_MUX_Subtract134_impl_0_parent_implementedSystem_port_2_cast <= SharedReg13_out;
   MUX_Subtract134_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg190_out_to_MUX_Subtract134_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg13_out_to_MUX_Subtract134_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract134_impl_0_out);

   Delay1No438_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract134_impl_0_out,
                 Y => Delay1No438_out);

SharedReg196_out_to_MUX_Subtract134_impl_1_parent_implementedSystem_port_1_cast <= SharedReg196_out;
SharedReg29_out_to_MUX_Subtract134_impl_1_parent_implementedSystem_port_2_cast <= SharedReg29_out;
   MUX_Subtract134_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg196_out_to_MUX_Subtract134_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg29_out_to_MUX_Subtract134_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract134_impl_1_out);

   Delay1No439_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract134_impl_1_out,
                 Y => Delay1No439_out);

Delay1No440_out_to_Subtract75_impl_parent_implementedSystem_port_0_cast <= Delay1No440_out;
Delay1No441_out_to_Subtract75_impl_parent_implementedSystem_port_1_cast <= Delay1No441_out;
   Subtract75_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract75_impl_out,
                 X => Delay1No440_out_to_Subtract75_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No441_out_to_Subtract75_impl_parent_implementedSystem_port_1_cast);

SharedReg207_out_to_MUX_Subtract75_impl_0_parent_implementedSystem_port_1_cast <= SharedReg207_out;
SharedReg14_out_to_MUX_Subtract75_impl_0_parent_implementedSystem_port_2_cast <= SharedReg14_out;
   MUX_Subtract75_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg207_out_to_MUX_Subtract75_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg14_out_to_MUX_Subtract75_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract75_impl_0_out);

   Delay1No440_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract75_impl_0_out,
                 Y => Delay1No440_out);

SharedReg213_out_to_MUX_Subtract75_impl_1_parent_implementedSystem_port_1_cast <= SharedReg213_out;
SharedReg30_out_to_MUX_Subtract75_impl_1_parent_implementedSystem_port_2_cast <= SharedReg30_out;
   MUX_Subtract75_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg213_out_to_MUX_Subtract75_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg30_out_to_MUX_Subtract75_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract75_impl_1_out);

   Delay1No441_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract75_impl_1_out,
                 Y => Delay1No441_out);

Delay1No442_out_to_Subtract135_impl_parent_implementedSystem_port_0_cast <= Delay1No442_out;
Delay1No443_out_to_Subtract135_impl_parent_implementedSystem_port_1_cast <= Delay1No443_out;
   Subtract135_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract135_impl_out,
                 X => Delay1No442_out_to_Subtract135_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No443_out_to_Subtract135_impl_parent_implementedSystem_port_1_cast);

SharedReg202_out_to_MUX_Subtract135_impl_0_parent_implementedSystem_port_1_cast <= SharedReg202_out;
SharedReg15_out_to_MUX_Subtract135_impl_0_parent_implementedSystem_port_2_cast <= SharedReg15_out;
   MUX_Subtract135_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg202_out_to_MUX_Subtract135_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg15_out_to_MUX_Subtract135_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract135_impl_0_out);

   Delay1No442_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract135_impl_0_out,
                 Y => Delay1No442_out);

SharedReg208_out_to_MUX_Subtract135_impl_1_parent_implementedSystem_port_1_cast <= SharedReg208_out;
SharedReg31_out_to_MUX_Subtract135_impl_1_parent_implementedSystem_port_2_cast <= SharedReg31_out;
   MUX_Subtract135_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg208_out_to_MUX_Subtract135_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg31_out_to_MUX_Subtract135_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract135_impl_1_out);

   Delay1No443_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract135_impl_1_out,
                 Y => Delay1No443_out);

Delay1No444_out_to_Subtract80_impl_parent_implementedSystem_port_0_cast <= Delay1No444_out;
Delay1No445_out_to_Subtract80_impl_parent_implementedSystem_port_1_cast <= Delay1No445_out;
   Subtract80_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract80_impl_out,
                 X => Delay1No444_out_to_Subtract80_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No445_out_to_Subtract80_impl_parent_implementedSystem_port_1_cast);

SharedReg81_out_to_MUX_Subtract80_impl_0_parent_implementedSystem_port_1_cast <= SharedReg81_out;
SharedReg83_out_to_MUX_Subtract80_impl_0_parent_implementedSystem_port_2_cast <= SharedReg83_out;
   MUX_Subtract80_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg81_out_to_MUX_Subtract80_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg83_out_to_MUX_Subtract80_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract80_impl_0_out);

   Delay1No444_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract80_impl_0_out,
                 Y => Delay1No444_out);

SharedReg165_out_to_MUX_Subtract80_impl_1_parent_implementedSystem_port_1_cast <= SharedReg165_out;
SharedReg214_out_to_MUX_Subtract80_impl_1_parent_implementedSystem_port_2_cast <= SharedReg214_out;
   MUX_Subtract80_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg165_out_to_MUX_Subtract80_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg214_out_to_MUX_Subtract80_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract80_impl_1_out);

   Delay1No445_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract80_impl_1_out,
                 Y => Delay1No445_out);

Delay1No446_out_to_Subtract140_impl_parent_implementedSystem_port_0_cast <= Delay1No446_out;
Delay1No447_out_to_Subtract140_impl_parent_implementedSystem_port_1_cast <= Delay1No447_out;
   Subtract140_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract140_impl_out,
                 X => Delay1No446_out_to_Subtract140_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No447_out_to_Subtract140_impl_parent_implementedSystem_port_1_cast);

SharedReg76_out_to_MUX_Subtract140_impl_0_parent_implementedSystem_port_1_cast <= SharedReg76_out;
SharedReg76_out_to_MUX_Subtract140_impl_0_parent_implementedSystem_port_2_cast <= SharedReg76_out;
   MUX_Subtract140_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg76_out_to_MUX_Subtract140_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg76_out_to_MUX_Subtract140_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract140_impl_0_out);

   Delay1No446_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract140_impl_0_out,
                 Y => Delay1No446_out);

SharedReg160_out_to_MUX_Subtract140_impl_1_parent_implementedSystem_port_1_cast <= SharedReg160_out;
SharedReg196_out_to_MUX_Subtract140_impl_1_parent_implementedSystem_port_2_cast <= SharedReg196_out;
   MUX_Subtract140_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg160_out_to_MUX_Subtract140_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg196_out_to_MUX_Subtract140_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => ModCount21_out,
                 oMux => MUX_Subtract140_impl_1_out);

   Delay1No447_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract140_impl_1_out,
                 Y => Delay1No447_out);
   Constant2_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant2_impl_out);
   Constant11_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant11_impl_out);
   Constant3_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant3_impl_out);
   Constant12_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant12_impl_out);
   Constant4_impl_instance: Constant_float_8_23_cosnpi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant4_impl_out);
   Constant13_impl_instance: Constant_float_8_23_sinnpi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant13_impl_out);
   Constant5_impl_instance: Constant_float_8_23_cosn3_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant5_impl_out);
   Constant14_impl_instance: Constant_float_8_23_sinn3_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant14_impl_out);
   Constant6_impl_instance: Constant_float_8_23_cosnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant6_impl_out);
   Constant15_impl_instance: Constant_float_8_23_sinnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant15_impl_out);
   Constant7_impl_instance: Constant_float_8_23_cosn5_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant7_impl_out);
   Constant16_impl_instance: Constant_float_8_23_sinn5_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant16_impl_out);
   Constant8_impl_instance: Constant_float_8_23_cosn3_mult_pi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant8_impl_out);
   Constant17_impl_instance: Constant_float_8_23_sinn3_mult_pi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant17_impl_out);
   Constant9_impl_instance: Constant_float_8_23_cosn7_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant9_impl_out);
   Constant18_impl_instance: Constant_float_8_23_sinn7_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant18_impl_out);
   Constant10_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant10_impl_out);
   Constant19_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant19_impl_out);
   Constant20_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant20_impl_out);
   Constant110_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant110_impl_out);
   Constant21_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant21_impl_out);
   Constant111_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant111_impl_out);
   Constant22_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant22_impl_out);
   Constant112_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant112_impl_out);
   Constant23_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant23_impl_out);
   Constant113_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant113_impl_out);
   Constant24_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant24_impl_out);
   Constant114_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant114_impl_out);
   Constant25_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant25_impl_out);
   Constant115_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant115_impl_out);
   Constant26_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant26_impl_out);
   Constant116_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant116_impl_out);
   Constant27_impl_instance: Constant_float_8_23_cosnpi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant27_impl_out);
   Constant117_impl_instance: Constant_float_8_23_sinnpi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant117_impl_out);
   Constant28_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant28_impl_out);
   Constant118_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant118_impl_out);
   Constant29_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant29_impl_out);
   Constant119_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant119_impl_out);
   Constant30_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant30_impl_out);
   Constant120_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant120_impl_out);
   Constant31_impl_instance: Constant_float_8_23_cosnpi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant31_impl_out);
   Constant121_impl_instance: Constant_float_8_23_sinnpi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant121_impl_out);
   Constant32_impl_instance: Constant_float_8_23_cosn3_mult_pi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant32_impl_out);
   Constant122_impl_instance: Constant_float_8_23_sinn3_mult_pi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant122_impl_out);
   Constant33_impl_instance: Constant_float_8_23_cosn3_mult_pi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant33_impl_out);
   Constant123_impl_instance: Constant_float_8_23_sinn3_mult_pi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant123_impl_out);
   Constant34_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant34_impl_out);
   Constant124_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant124_impl_out);
   Constant35_impl_instance: Constant_float_8_23_cosnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant35_impl_out);
   Constant125_impl_instance: Constant_float_8_23_sinnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant125_impl_out);
   Constant36_impl_instance: Constant_float_8_23_cosnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant36_impl_out);
   Constant126_impl_instance: Constant_float_8_23_sinnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant126_impl_out);
   Constant37_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant37_impl_out);
   Constant127_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant127_impl_out);
   Constant38_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant38_impl_out);
   Constant128_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant128_impl_out);
   Constant39_impl_instance: Constant_float_8_23_cosnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant39_impl_out);
   Constant129_impl_instance: Constant_float_8_23_sinnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant129_impl_out);
   Constant40_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant40_impl_out);
   Constant130_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant130_impl_out);
   Constant41_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant41_impl_out);
   Constant131_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant131_impl_out);
   Constant42_impl_instance: Constant_float_8_23_cosnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant42_impl_out);
   Constant132_impl_instance: Constant_float_8_23_sinnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant132_impl_out);
   Constant43_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant43_impl_out);
   Constant133_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant133_impl_out);
   Constant44_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant44_impl_out);
   Constant134_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant134_impl_out);
   Constant45_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant45_impl_out);
   Constant135_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant135_impl_out);
   Constant46_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant46_impl_out);
   Constant136_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant136_impl_out);
   Constant47_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant47_impl_out);
   Constant137_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant137_impl_out);
   Constant48_impl_instance: Constant_float_8_23_cosnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant48_impl_out);
   Constant138_impl_instance: Constant_float_8_23_sinnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant138_impl_out);
   Constant49_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant49_impl_out);
   Constant139_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant139_impl_out);
   Constant50_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant50_impl_out);
   Constant140_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant140_impl_out);
   Constant51_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant51_impl_out);
   Constant141_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant141_impl_out);
   Constant52_impl_instance: Constant_float_8_23_cosnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant52_impl_out);
   Constant142_impl_instance: Constant_float_8_23_sinnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant142_impl_out);
   Constant53_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant53_impl_out);
   Constant143_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant143_impl_out);
   Constant54_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant54_impl_out);
   Constant144_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant144_impl_out);
   Constant55_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant55_impl_out);
   Constant145_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant145_impl_out);
   Constant56_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant56_impl_out);
   Constant146_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant146_impl_out);
   Constant57_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant57_impl_out);
   Constant147_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant147_impl_out);
   Constant_impl_instance: Constant_float_8_23_cosnpi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant_impl_out);
   Constant1_impl_instance: Constant_float_8_23_sinnpi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant1_impl_out);

   Delay2No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg_out,
                 Y => Delay2No_out);

   Delay2No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1_out,
                 Y => Delay2No1_out);

   Delay2No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg4_out,
                 Y => Delay2No2_out);

   Delay2No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg5_out,
                 Y => Delay2No3_out);

   Delay2No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg8_out,
                 Y => Delay2No4_out);

   Delay2No5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg9_out,
                 Y => Delay2No5_out);

   Delay2No6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg12_out,
                 Y => Delay2No6_out);

   Delay2No7_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg13_out,
                 Y => Delay2No7_out);

   Delay2No8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg16_out,
                 Y => Delay2No8_out);

   Delay2No9_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg17_out,
                 Y => Delay2No9_out);

   Delay2No10_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg20_out,
                 Y => Delay2No10_out);

   Delay2No11_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg21_out,
                 Y => Delay2No11_out);

   Delay2No12_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg24_out,
                 Y => Delay2No12_out);

   Delay2No13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg25_out,
                 Y => Delay2No13_out);

   Delay2No14_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg28_out,
                 Y => Delay2No14_out);

   Delay2No15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg29_out,
                 Y => Delay2No15_out);

   Delay2No40_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg130_out,
                 Y => Delay2No40_out);

   Delay2No41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg135_out,
                 Y => Delay2No41_out);

   Delay2No42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg142_out,
                 Y => Delay2No42_out);

   Delay2No43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg147_out,
                 Y => Delay2No43_out);

   Delay2No44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg148_out,
                 Y => Delay2No44_out);

   Delay2No45_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg153_out,
                 Y => Delay2No45_out);

   Delay2No46_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg154_out,
                 Y => Delay2No46_out);

   Delay2No47_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg159_out,
                 Y => Delay2No47_out);

   Delay2No48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg166_out,
                 Y => Delay2No48_out);

   Delay2No49_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg171_out,
                 Y => Delay2No49_out);

   Delay2No50_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg172_out,
                 Y => Delay2No50_out);

   Delay2No51_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg177_out,
                 Y => Delay2No51_out);

   Delay2No52_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg184_out,
                 Y => Delay2No52_out);

   Delay2No53_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg189_out,
                 Y => Delay2No53_out);

   Delay2No54_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg190_out,
                 Y => Delay2No54_out);

   Delay2No55_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg195_out,
                 Y => Delay2No55_out);

   SharedReg_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x0_re_out,
                 Y => SharedReg_out);

   SharedReg1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x0_im_out,
                 Y => SharedReg1_out);

   SharedReg2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x1_re_out,
                 Y => SharedReg2_out);

   SharedReg3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x1_im_out,
                 Y => SharedReg3_out);

   SharedReg4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x2_re_out,
                 Y => SharedReg4_out);

   SharedReg5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x2_im_out,
                 Y => SharedReg5_out);

   SharedReg6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x3_re_out,
                 Y => SharedReg6_out);

   SharedReg7_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x3_im_out,
                 Y => SharedReg7_out);

   SharedReg8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x4_re_out,
                 Y => SharedReg8_out);

   SharedReg9_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x4_im_out,
                 Y => SharedReg9_out);

   SharedReg10_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x5_re_out,
                 Y => SharedReg10_out);

   SharedReg11_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x5_im_out,
                 Y => SharedReg11_out);

   SharedReg12_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x6_re_out,
                 Y => SharedReg12_out);

   SharedReg13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x6_im_out,
                 Y => SharedReg13_out);

   SharedReg14_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x7_re_out,
                 Y => SharedReg14_out);

   SharedReg15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x7_im_out,
                 Y => SharedReg15_out);

   SharedReg16_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x8_re_out,
                 Y => SharedReg16_out);

   SharedReg17_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x8_im_out,
                 Y => SharedReg17_out);

   SharedReg18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x9_re_out,
                 Y => SharedReg18_out);

   SharedReg19_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x9_im_out,
                 Y => SharedReg19_out);

   SharedReg20_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x10_re_out,
                 Y => SharedReg20_out);

   SharedReg21_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x10_im_out,
                 Y => SharedReg21_out);

   SharedReg22_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x11_re_out,
                 Y => SharedReg22_out);

   SharedReg23_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x11_im_out,
                 Y => SharedReg23_out);

   SharedReg24_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x12_re_out,
                 Y => SharedReg24_out);

   SharedReg25_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x12_im_out,
                 Y => SharedReg25_out);

   SharedReg26_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x13_re_out,
                 Y => SharedReg26_out);

   SharedReg27_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x13_im_out,
                 Y => SharedReg27_out);

   SharedReg28_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x14_re_out,
                 Y => SharedReg28_out);

   SharedReg29_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x14_im_out,
                 Y => SharedReg29_out);

   SharedReg30_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x15_re_out,
                 Y => SharedReg30_out);

   SharedReg31_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x15_im_out,
                 Y => SharedReg31_out);

   SharedReg32_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_impl_out,
                 Y => SharedReg32_out);

   SharedReg33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_impl_out,
                 Y => SharedReg33_out);

   SharedReg34_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add12_impl_out,
                 Y => SharedReg34_out);

   SharedReg35_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add13_impl_out,
                 Y => SharedReg35_out);

   SharedReg36_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add14_impl_out,
                 Y => SharedReg36_out);

   SharedReg37_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add6_impl_out,
                 Y => SharedReg37_out);

   SharedReg38_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add15_impl_out,
                 Y => SharedReg38_out);

   SharedReg39_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add7_impl_out,
                 Y => SharedReg39_out);

   SharedReg40_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add16_impl_out,
                 Y => SharedReg40_out);

   SharedReg41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add8_impl_out,
                 Y => SharedReg41_out);

   SharedReg42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add9_impl_out,
                 Y => SharedReg42_out);

   SharedReg43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add18_impl_out,
                 Y => SharedReg43_out);

   SharedReg44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add20_impl_out,
                 Y => SharedReg44_out);

   SharedReg45_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg44_out,
                 Y => SharedReg45_out);

   SharedReg46_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add110_impl_out,
                 Y => SharedReg46_out);

   SharedReg47_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg46_out,
                 Y => SharedReg47_out);

   SharedReg48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add22_impl_out,
                 Y => SharedReg48_out);

   SharedReg49_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg48_out,
                 Y => SharedReg49_out);

   SharedReg50_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add112_impl_out,
                 Y => SharedReg50_out);

   SharedReg51_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg50_out,
                 Y => SharedReg51_out);

   SharedReg52_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add24_impl_out,
                 Y => SharedReg52_out);

   SharedReg53_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg52_out,
                 Y => SharedReg53_out);

   SharedReg54_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add114_impl_out,
                 Y => SharedReg54_out);

   SharedReg55_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg54_out,
                 Y => SharedReg55_out);

   SharedReg56_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add25_impl_out,
                 Y => SharedReg56_out);

   SharedReg57_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg56_out,
                 Y => SharedReg57_out);

   SharedReg58_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add115_impl_out,
                 Y => SharedReg58_out);

   SharedReg59_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg58_out,
                 Y => SharedReg59_out);

   SharedReg60_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add26_impl_out,
                 Y => SharedReg60_out);

   SharedReg61_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg60_out,
                 Y => SharedReg61_out);

   SharedReg62_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add116_impl_out,
                 Y => SharedReg62_out);

   SharedReg63_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg62_out,
                 Y => SharedReg63_out);

   SharedReg64_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add27_impl_out,
                 Y => SharedReg64_out);

   SharedReg65_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg64_out,
                 Y => SharedReg65_out);

   SharedReg66_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add117_impl_out,
                 Y => SharedReg66_out);

   SharedReg67_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg66_out,
                 Y => SharedReg67_out);

   SharedReg68_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add34_impl_out,
                 Y => SharedReg68_out);

   SharedReg69_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add124_impl_out,
                 Y => SharedReg69_out);

   SharedReg70_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add126_impl_out,
                 Y => SharedReg70_out);

   SharedReg71_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add37_impl_out,
                 Y => SharedReg71_out);

   SharedReg72_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add127_impl_out,
                 Y => SharedReg72_out);

   SharedReg73_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add129_impl_out,
                 Y => SharedReg73_out);

   SharedReg74_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add41_impl_out,
                 Y => SharedReg74_out);

   SharedReg75_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add131_impl_out,
                 Y => SharedReg75_out);

   SharedReg76_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add43_impl_out,
                 Y => SharedReg76_out);

   SharedReg77_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_impl_out,
                 Y => SharedReg77_out);

   SharedReg78_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product11_impl_out,
                 Y => SharedReg78_out);

   SharedReg79_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_impl_out,
                 Y => SharedReg79_out);

   SharedReg80_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product31_impl_out,
                 Y => SharedReg80_out);

   SharedReg81_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_impl_out,
                 Y => SharedReg81_out);

   SharedReg82_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_impl_out,
                 Y => SharedReg82_out);

   SharedReg83_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract3_impl_out,
                 Y => SharedReg83_out);

   SharedReg84_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add45_impl_out,
                 Y => SharedReg84_out);

   SharedReg85_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product6_impl_out,
                 Y => SharedReg85_out);

   SharedReg86_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product13_impl_out,
                 Y => SharedReg86_out);

   SharedReg87_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product23_impl_out,
                 Y => SharedReg87_out);

   SharedReg88_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product33_impl_out,
                 Y => SharedReg88_out);

   SharedReg89_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract4_impl_out,
                 Y => SharedReg89_out);

   SharedReg90_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add46_impl_out,
                 Y => SharedReg90_out);

   SharedReg91_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product7_impl_out,
                 Y => SharedReg91_out);

   SharedReg92_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product14_impl_out,
                 Y => SharedReg92_out);

   SharedReg93_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product24_impl_out,
                 Y => SharedReg93_out);

   SharedReg94_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add47_impl_out,
                 Y => SharedReg94_out);

   SharedReg95_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product8_impl_out,
                 Y => SharedReg95_out);

   SharedReg96_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product15_impl_out,
                 Y => SharedReg96_out);

   SharedReg97_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product25_impl_out,
                 Y => SharedReg97_out);

   SharedReg98_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product35_impl_out,
                 Y => SharedReg98_out);

   SharedReg99_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract6_impl_out,
                 Y => SharedReg99_out);

   SharedReg100_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add48_impl_out,
                 Y => SharedReg100_out);

   SharedReg101_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product9_impl_out,
                 Y => SharedReg101_out);

   SharedReg102_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product16_impl_out,
                 Y => SharedReg102_out);

   SharedReg103_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product26_impl_out,
                 Y => SharedReg103_out);

   SharedReg104_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product36_impl_out,
                 Y => SharedReg104_out);

   SharedReg105_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract7_impl_out,
                 Y => SharedReg105_out);

   SharedReg106_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add49_impl_out,
                 Y => SharedReg106_out);

   SharedReg107_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product10_impl_out,
                 Y => SharedReg107_out);

   SharedReg108_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product17_impl_out,
                 Y => SharedReg108_out);

   SharedReg109_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product27_impl_out,
                 Y => SharedReg109_out);

   SharedReg110_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product37_impl_out,
                 Y => SharedReg110_out);

   SharedReg111_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract8_impl_out,
                 Y => SharedReg111_out);

   SharedReg112_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add50_impl_out,
                 Y => SharedReg112_out);

   SharedReg113_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product18_impl_out,
                 Y => SharedReg113_out);

   SharedReg114_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product19_impl_out,
                 Y => SharedReg114_out);

   SharedReg115_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product28_impl_out,
                 Y => SharedReg115_out);

   SharedReg116_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product38_impl_out,
                 Y => SharedReg116_out);

   SharedReg117_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract9_impl_out,
                 Y => SharedReg117_out);

   SharedReg118_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add52_impl_out,
                 Y => SharedReg118_out);

   SharedReg119_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product30_impl_out,
                 Y => SharedReg119_out);

   SharedReg120_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product111_impl_out,
                 Y => SharedReg120_out);

   SharedReg121_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product210_impl_out,
                 Y => SharedReg121_out);

   SharedReg122_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product310_impl_out,
                 Y => SharedReg122_out);

   SharedReg123_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract11_impl_out,
                 Y => SharedReg123_out);

   SharedReg124_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add53_impl_out,
                 Y => SharedReg124_out);

   SharedReg125_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product40_impl_out,
                 Y => SharedReg125_out);

   SharedReg126_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product112_impl_out,
                 Y => SharedReg126_out);

   SharedReg127_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product211_impl_out,
                 Y => SharedReg127_out);

   SharedReg128_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product311_impl_out,
                 Y => SharedReg128_out);

   SharedReg129_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract12_impl_out,
                 Y => SharedReg129_out);

   SharedReg130_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add54_impl_out,
                 Y => SharedReg130_out);

   SharedReg131_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product41_impl_out,
                 Y => SharedReg131_out);

   SharedReg132_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product113_impl_out,
                 Y => SharedReg132_out);

   SharedReg133_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product212_impl_out,
                 Y => SharedReg133_out);

   SharedReg134_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product312_impl_out,
                 Y => SharedReg134_out);

   SharedReg135_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract13_impl_out,
                 Y => SharedReg135_out);

   SharedReg136_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add56_impl_out,
                 Y => SharedReg136_out);

   SharedReg137_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product43_impl_out,
                 Y => SharedReg137_out);

   SharedReg138_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product115_impl_out,
                 Y => SharedReg138_out);

   SharedReg139_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product214_impl_out,
                 Y => SharedReg139_out);

   SharedReg140_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product314_impl_out,
                 Y => SharedReg140_out);

   SharedReg141_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract15_impl_out,
                 Y => SharedReg141_out);

   SharedReg142_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add57_impl_out,
                 Y => SharedReg142_out);

   SharedReg143_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product44_impl_out,
                 Y => SharedReg143_out);

   SharedReg144_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product116_impl_out,
                 Y => SharedReg144_out);

   SharedReg145_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product215_impl_out,
                 Y => SharedReg145_out);

   SharedReg146_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product315_impl_out,
                 Y => SharedReg146_out);

   SharedReg147_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract16_impl_out,
                 Y => SharedReg147_out);

   SharedReg148_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add58_impl_out,
                 Y => SharedReg148_out);

   SharedReg149_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product45_impl_out,
                 Y => SharedReg149_out);

   SharedReg150_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product117_impl_out,
                 Y => SharedReg150_out);

   SharedReg151_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product216_impl_out,
                 Y => SharedReg151_out);

   SharedReg152_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product316_impl_out,
                 Y => SharedReg152_out);

   SharedReg153_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract17_impl_out,
                 Y => SharedReg153_out);

   SharedReg154_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add59_impl_out,
                 Y => SharedReg154_out);

   SharedReg155_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product46_impl_out,
                 Y => SharedReg155_out);

   SharedReg156_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product118_impl_out,
                 Y => SharedReg156_out);

   SharedReg157_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product217_impl_out,
                 Y => SharedReg157_out);

   SharedReg158_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product317_impl_out,
                 Y => SharedReg158_out);

   SharedReg159_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract18_impl_out,
                 Y => SharedReg159_out);

   SharedReg160_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add61_impl_out,
                 Y => SharedReg160_out);

   SharedReg161_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product48_impl_out,
                 Y => SharedReg161_out);

   SharedReg162_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product120_impl_out,
                 Y => SharedReg162_out);

   SharedReg163_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product219_impl_out,
                 Y => SharedReg163_out);

   SharedReg164_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product319_impl_out,
                 Y => SharedReg164_out);

   SharedReg165_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract20_impl_out,
                 Y => SharedReg165_out);

   SharedReg166_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add63_impl_out,
                 Y => SharedReg166_out);

   SharedReg167_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product50_impl_out,
                 Y => SharedReg167_out);

   SharedReg168_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product122_impl_out,
                 Y => SharedReg168_out);

   SharedReg169_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product221_impl_out,
                 Y => SharedReg169_out);

   SharedReg170_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product321_impl_out,
                 Y => SharedReg170_out);

   SharedReg171_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract22_impl_out,
                 Y => SharedReg171_out);

   SharedReg172_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add65_impl_out,
                 Y => SharedReg172_out);

   SharedReg173_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product52_impl_out,
                 Y => SharedReg173_out);

   SharedReg174_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product124_impl_out,
                 Y => SharedReg174_out);

   SharedReg175_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product223_impl_out,
                 Y => SharedReg175_out);

   SharedReg176_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product323_impl_out,
                 Y => SharedReg176_out);

   SharedReg177_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract24_impl_out,
                 Y => SharedReg177_out);

   SharedReg178_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add66_impl_out,
                 Y => SharedReg178_out);

   SharedReg179_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product53_impl_out,
                 Y => SharedReg179_out);

   SharedReg180_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product125_impl_out,
                 Y => SharedReg180_out);

   SharedReg181_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product224_impl_out,
                 Y => SharedReg181_out);

   SharedReg182_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product324_impl_out,
                 Y => SharedReg182_out);

   SharedReg183_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract25_impl_out,
                 Y => SharedReg183_out);

   SharedReg184_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add67_impl_out,
                 Y => SharedReg184_out);

   SharedReg185_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product54_impl_out,
                 Y => SharedReg185_out);

   SharedReg186_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product126_impl_out,
                 Y => SharedReg186_out);

   SharedReg187_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product225_impl_out,
                 Y => SharedReg187_out);

   SharedReg188_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product325_impl_out,
                 Y => SharedReg188_out);

   SharedReg189_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract26_impl_out,
                 Y => SharedReg189_out);

   SharedReg190_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add68_impl_out,
                 Y => SharedReg190_out);

   SharedReg191_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product55_impl_out,
                 Y => SharedReg191_out);

   SharedReg192_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product127_impl_out,
                 Y => SharedReg192_out);

   SharedReg193_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product226_impl_out,
                 Y => SharedReg193_out);

   SharedReg194_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product326_impl_out,
                 Y => SharedReg194_out);

   SharedReg195_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract27_impl_out,
                 Y => SharedReg195_out);

   SharedReg196_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add83_impl_out,
                 Y => SharedReg196_out);

   SharedReg197_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product70_impl_out,
                 Y => SharedReg197_out);

   SharedReg198_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product142_impl_out,
                 Y => SharedReg198_out);

   SharedReg199_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product241_impl_out,
                 Y => SharedReg199_out);

   SharedReg200_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product341_impl_out,
                 Y => SharedReg200_out);

   SharedReg201_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract42_impl_out,
                 Y => SharedReg201_out);

   SharedReg202_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add84_impl_out,
                 Y => SharedReg202_out);

   SharedReg203_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product71_impl_out,
                 Y => SharedReg203_out);

   SharedReg204_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product143_impl_out,
                 Y => SharedReg204_out);

   SharedReg205_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product242_impl_out,
                 Y => SharedReg205_out);

   SharedReg206_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product342_impl_out,
                 Y => SharedReg206_out);

   SharedReg207_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract43_impl_out,
                 Y => SharedReg207_out);

   SharedReg208_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add85_impl_out,
                 Y => SharedReg208_out);

   SharedReg209_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product72_impl_out,
                 Y => SharedReg209_out);

   SharedReg210_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product144_impl_out,
                 Y => SharedReg210_out);

   SharedReg211_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product243_impl_out,
                 Y => SharedReg211_out);

   SharedReg212_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product343_impl_out,
                 Y => SharedReg212_out);

   SharedReg213_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract44_impl_out,
                 Y => SharedReg213_out);

   SharedReg214_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract45_impl_out,
                 Y => SharedReg214_out);

   SharedReg215_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add87_impl_out,
                 Y => SharedReg215_out);

   SharedReg216_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product74_impl_out,
                 Y => SharedReg216_out);

   SharedReg217_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product146_impl_out,
                 Y => SharedReg217_out);

   SharedReg218_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product245_impl_out,
                 Y => SharedReg218_out);

   SharedReg219_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product345_impl_out,
                 Y => SharedReg219_out);

   SharedReg220_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract46_impl_out,
                 Y => SharedReg220_out);

   SharedReg221_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract47_impl_out,
                 Y => SharedReg221_out);

   SharedReg222_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract48_impl_out,
                 Y => SharedReg222_out);

   SharedReg223_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract49_impl_out,
                 Y => SharedReg223_out);

   SharedReg224_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract50_impl_out,
                 Y => SharedReg224_out);

   SharedReg225_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract52_impl_out,
                 Y => SharedReg225_out);

   SharedReg226_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract112_impl_out,
                 Y => SharedReg226_out);

   SharedReg227_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract114_impl_out,
                 Y => SharedReg227_out);

   SharedReg228_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract55_impl_out,
                 Y => SharedReg228_out);

   SharedReg229_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract115_impl_out,
                 Y => SharedReg229_out);

   SharedReg230_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract56_impl_out,
                 Y => SharedReg230_out);

   SharedReg231_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract116_impl_out,
                 Y => SharedReg231_out);

   SharedReg232_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract57_impl_out,
                 Y => SharedReg232_out);

   SharedReg233_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract117_impl_out,
                 Y => SharedReg233_out);

   SharedReg234_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract59_impl_out,
                 Y => SharedReg234_out);

   SharedReg235_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg234_out,
                 Y => SharedReg235_out);

   SharedReg236_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract119_impl_out,
                 Y => SharedReg236_out);

   SharedReg237_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg236_out,
                 Y => SharedReg237_out);

   SharedReg238_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract62_impl_out,
                 Y => SharedReg238_out);

   SharedReg239_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract122_impl_out,
                 Y => SharedReg239_out);

   SharedReg240_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract63_impl_out,
                 Y => SharedReg240_out);

   SharedReg241_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg240_out,
                 Y => SharedReg241_out);

   SharedReg242_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract123_impl_out,
                 Y => SharedReg242_out);

   SharedReg243_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg242_out,
                 Y => SharedReg243_out);

   SharedReg244_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract127_impl_out,
                 Y => SharedReg244_out);

   SharedReg245_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract68_impl_out,
                 Y => SharedReg245_out);

   SharedReg246_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract71_impl_out,
                 Y => SharedReg246_out);

   SharedReg247_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract131_impl_out,
                 Y => SharedReg247_out);

   SharedReg248_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract72_impl_out,
                 Y => SharedReg248_out);

   SharedReg249_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract132_impl_out,
                 Y => SharedReg249_out);

   SharedReg250_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract74_impl_out,
                 Y => SharedReg250_out);

   SharedReg251_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract134_impl_out,
                 Y => SharedReg251_out);

   SharedReg252_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract75_impl_out,
                 Y => SharedReg252_out);

   SharedReg253_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract135_impl_out,
                 Y => SharedReg253_out);

   SharedReg254_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract80_impl_out,
                 Y => SharedReg254_out);

   SharedReg255_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract140_impl_out,
                 Y => SharedReg255_out);

   SharedReg256_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant2_impl_out,
                 Y => SharedReg256_out);

   SharedReg257_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant11_impl_out,
                 Y => SharedReg257_out);

   SharedReg258_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant3_impl_out,
                 Y => SharedReg258_out);

   SharedReg259_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant12_impl_out,
                 Y => SharedReg259_out);

   SharedReg260_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant4_impl_out,
                 Y => SharedReg260_out);

   SharedReg261_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant13_impl_out,
                 Y => SharedReg261_out);

   SharedReg262_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant5_impl_out,
                 Y => SharedReg262_out);

   SharedReg263_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant14_impl_out,
                 Y => SharedReg263_out);

   SharedReg264_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant6_impl_out,
                 Y => SharedReg264_out);

   SharedReg265_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant15_impl_out,
                 Y => SharedReg265_out);

   SharedReg266_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant7_impl_out,
                 Y => SharedReg266_out);

   SharedReg267_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant16_impl_out,
                 Y => SharedReg267_out);

   SharedReg268_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant8_impl_out,
                 Y => SharedReg268_out);

   SharedReg269_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant17_impl_out,
                 Y => SharedReg269_out);

   SharedReg270_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant9_impl_out,
                 Y => SharedReg270_out);

   SharedReg271_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant18_impl_out,
                 Y => SharedReg271_out);

   SharedReg272_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant10_impl_out,
                 Y => SharedReg272_out);

   SharedReg273_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant19_impl_out,
                 Y => SharedReg273_out);

   SharedReg274_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant20_impl_out,
                 Y => SharedReg274_out);

   SharedReg275_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant110_impl_out,
                 Y => SharedReg275_out);

   SharedReg276_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant21_impl_out,
                 Y => SharedReg276_out);

   SharedReg277_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant111_impl_out,
                 Y => SharedReg277_out);

   SharedReg278_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant22_impl_out,
                 Y => SharedReg278_out);

   SharedReg279_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant112_impl_out,
                 Y => SharedReg279_out);

   SharedReg280_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant23_impl_out,
                 Y => SharedReg280_out);

   SharedReg281_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant113_impl_out,
                 Y => SharedReg281_out);

   SharedReg282_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant24_impl_out,
                 Y => SharedReg282_out);

   SharedReg283_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant114_impl_out,
                 Y => SharedReg283_out);

   SharedReg284_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant25_impl_out,
                 Y => SharedReg284_out);

   SharedReg285_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant115_impl_out,
                 Y => SharedReg285_out);

   SharedReg286_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant26_impl_out,
                 Y => SharedReg286_out);

   SharedReg287_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant116_impl_out,
                 Y => SharedReg287_out);

   SharedReg288_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant27_impl_out,
                 Y => SharedReg288_out);

   SharedReg289_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant117_impl_out,
                 Y => SharedReg289_out);

   SharedReg290_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant28_impl_out,
                 Y => SharedReg290_out);

   SharedReg291_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant118_impl_out,
                 Y => SharedReg291_out);

   SharedReg292_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant29_impl_out,
                 Y => SharedReg292_out);

   SharedReg293_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant119_impl_out,
                 Y => SharedReg293_out);

   SharedReg294_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant30_impl_out,
                 Y => SharedReg294_out);

   SharedReg295_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant120_impl_out,
                 Y => SharedReg295_out);

   SharedReg296_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant31_impl_out,
                 Y => SharedReg296_out);

   SharedReg297_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant121_impl_out,
                 Y => SharedReg297_out);

   SharedReg298_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant32_impl_out,
                 Y => SharedReg298_out);

   SharedReg299_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant122_impl_out,
                 Y => SharedReg299_out);

   SharedReg300_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant33_impl_out,
                 Y => SharedReg300_out);

   SharedReg301_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant123_impl_out,
                 Y => SharedReg301_out);

   SharedReg302_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant34_impl_out,
                 Y => SharedReg302_out);

   SharedReg303_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant124_impl_out,
                 Y => SharedReg303_out);

   SharedReg304_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant35_impl_out,
                 Y => SharedReg304_out);

   SharedReg305_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant125_impl_out,
                 Y => SharedReg305_out);

   SharedReg306_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant36_impl_out,
                 Y => SharedReg306_out);

   SharedReg307_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant126_impl_out,
                 Y => SharedReg307_out);

   SharedReg308_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant37_impl_out,
                 Y => SharedReg308_out);

   SharedReg309_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant127_impl_out,
                 Y => SharedReg309_out);

   SharedReg310_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant38_impl_out,
                 Y => SharedReg310_out);

   SharedReg311_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant128_impl_out,
                 Y => SharedReg311_out);

   SharedReg312_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant39_impl_out,
                 Y => SharedReg312_out);

   SharedReg313_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant129_impl_out,
                 Y => SharedReg313_out);

   SharedReg314_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant40_impl_out,
                 Y => SharedReg314_out);

   SharedReg315_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant130_impl_out,
                 Y => SharedReg315_out);

   SharedReg316_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant41_impl_out,
                 Y => SharedReg316_out);

   SharedReg317_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant131_impl_out,
                 Y => SharedReg317_out);

   SharedReg318_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant42_impl_out,
                 Y => SharedReg318_out);

   SharedReg319_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant132_impl_out,
                 Y => SharedReg319_out);

   SharedReg320_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant43_impl_out,
                 Y => SharedReg320_out);

   SharedReg321_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant133_impl_out,
                 Y => SharedReg321_out);

   SharedReg322_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant44_impl_out,
                 Y => SharedReg322_out);

   SharedReg323_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant134_impl_out,
                 Y => SharedReg323_out);

   SharedReg324_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant45_impl_out,
                 Y => SharedReg324_out);

   SharedReg325_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant135_impl_out,
                 Y => SharedReg325_out);

   SharedReg326_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant46_impl_out,
                 Y => SharedReg326_out);

   SharedReg327_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant136_impl_out,
                 Y => SharedReg327_out);

   SharedReg328_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant47_impl_out,
                 Y => SharedReg328_out);

   SharedReg329_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant137_impl_out,
                 Y => SharedReg329_out);

   SharedReg330_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant48_impl_out,
                 Y => SharedReg330_out);

   SharedReg331_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant138_impl_out,
                 Y => SharedReg331_out);

   SharedReg332_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant49_impl_out,
                 Y => SharedReg332_out);

   SharedReg333_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant139_impl_out,
                 Y => SharedReg333_out);

   SharedReg334_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant50_impl_out,
                 Y => SharedReg334_out);

   SharedReg335_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant140_impl_out,
                 Y => SharedReg335_out);

   SharedReg336_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant51_impl_out,
                 Y => SharedReg336_out);

   SharedReg337_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant141_impl_out,
                 Y => SharedReg337_out);

   SharedReg338_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant52_impl_out,
                 Y => SharedReg338_out);

   SharedReg339_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant142_impl_out,
                 Y => SharedReg339_out);

   SharedReg340_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant53_impl_out,
                 Y => SharedReg340_out);

   SharedReg341_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant143_impl_out,
                 Y => SharedReg341_out);

   SharedReg342_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant54_impl_out,
                 Y => SharedReg342_out);

   SharedReg343_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant144_impl_out,
                 Y => SharedReg343_out);

   SharedReg344_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant55_impl_out,
                 Y => SharedReg344_out);

   SharedReg345_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant145_impl_out,
                 Y => SharedReg345_out);

   SharedReg346_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant56_impl_out,
                 Y => SharedReg346_out);

   SharedReg347_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant146_impl_out,
                 Y => SharedReg347_out);

   SharedReg348_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant57_impl_out,
                 Y => SharedReg348_out);

   SharedReg349_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant147_impl_out,
                 Y => SharedReg349_out);

   SharedReg350_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant_impl_out,
                 Y => SharedReg350_out);

   SharedReg351_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant1_impl_out,
                 Y => SharedReg351_out);
end architecture;



library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity implementedSystem_toplevel_wrapper is
  port (
    clk, rst : in std_logic;
    shared_input : in std_logic_vector(31 downto 0);
    x0_re_enable : in std_logic;
    x0_im_enable : in std_logic;
    x1_re_enable : in std_logic;
    x1_im_enable : in std_logic;
    x2_re_enable : in std_logic;
    x2_im_enable : in std_logic;
    x3_re_enable : in std_logic;
    x3_im_enable : in std_logic;
    x4_re_enable : in std_logic;
    x4_im_enable : in std_logic;
    x5_re_enable : in std_logic;
    x5_im_enable : in std_logic;
    x6_re_enable : in std_logic;
    x6_im_enable : in std_logic;
    x7_re_enable : in std_logic;
    x7_im_enable : in std_logic;
    x8_re_enable : in std_logic;
    x8_im_enable : in std_logic;
    x9_re_enable : in std_logic;
    x9_im_enable : in std_logic;
    x10_re_enable : in std_logic;
    x10_im_enable : in std_logic;
    x11_re_enable : in std_logic;
    x11_im_enable : in std_logic;
    x12_re_enable : in std_logic;
    x12_im_enable : in std_logic;
    x13_re_enable : in std_logic;
    x13_im_enable : in std_logic;
    x14_re_enable : in std_logic;
    x14_im_enable : in std_logic;
    x15_re_enable : in std_logic;
    x15_im_enable : in std_logic;
    output_select : in std_logic_vector(4 downto 0);
    shared_output : out std_logic_vector(31 downto 0)
  );
end entity;

architecture implementedSystem_toplevel_wrapper of implementedSystem_toplevel_wrapper is
  signal x0_re_DUT_in : std_logic_vector(31 downto 0);
  signal x0_im_DUT_in : std_logic_vector(31 downto 0);
  signal x1_re_DUT_in : std_logic_vector(31 downto 0);
  signal x1_im_DUT_in : std_logic_vector(31 downto 0);
  signal x2_re_DUT_in : std_logic_vector(31 downto 0);
  signal x2_im_DUT_in : std_logic_vector(31 downto 0);
  signal x3_re_DUT_in : std_logic_vector(31 downto 0);
  signal x3_im_DUT_in : std_logic_vector(31 downto 0);
  signal x4_re_DUT_in : std_logic_vector(31 downto 0);
  signal x4_im_DUT_in : std_logic_vector(31 downto 0);
  signal x5_re_DUT_in : std_logic_vector(31 downto 0);
  signal x5_im_DUT_in : std_logic_vector(31 downto 0);
  signal x6_re_DUT_in : std_logic_vector(31 downto 0);
  signal x6_im_DUT_in : std_logic_vector(31 downto 0);
  signal x7_re_DUT_in : std_logic_vector(31 downto 0);
  signal x7_im_DUT_in : std_logic_vector(31 downto 0);
  signal x8_re_DUT_in : std_logic_vector(31 downto 0);
  signal x8_im_DUT_in : std_logic_vector(31 downto 0);
  signal x9_re_DUT_in : std_logic_vector(31 downto 0);
  signal x9_im_DUT_in : std_logic_vector(31 downto 0);
  signal x10_re_DUT_in : std_logic_vector(31 downto 0);
  signal x10_im_DUT_in : std_logic_vector(31 downto 0);
  signal x11_re_DUT_in : std_logic_vector(31 downto 0);
  signal x11_im_DUT_in : std_logic_vector(31 downto 0);
  signal x12_re_DUT_in : std_logic_vector(31 downto 0);
  signal x12_im_DUT_in : std_logic_vector(31 downto 0);
  signal x13_re_DUT_in : std_logic_vector(31 downto 0);
  signal x13_im_DUT_in : std_logic_vector(31 downto 0);
  signal x14_re_DUT_in : std_logic_vector(31 downto 0);
  signal x14_im_DUT_in : std_logic_vector(31 downto 0);
  signal x15_re_DUT_in : std_logic_vector(31 downto 0);
  signal x15_im_DUT_in : std_logic_vector(31 downto 0);
  signal y0_re_DUT_out : std_logic_vector(31 downto 0);
  signal y0_im_DUT_out : std_logic_vector(31 downto 0);
  signal y1_re_DUT_out : std_logic_vector(31 downto 0);
  signal y1_im_DUT_out : std_logic_vector(31 downto 0);
  signal y2_re_DUT_out : std_logic_vector(31 downto 0);
  signal y2_im_DUT_out : std_logic_vector(31 downto 0);
  signal y3_re_DUT_out : std_logic_vector(31 downto 0);
  signal y3_im_DUT_out : std_logic_vector(31 downto 0);
  signal y4_re_DUT_out : std_logic_vector(31 downto 0);
  signal y4_im_DUT_out : std_logic_vector(31 downto 0);
  signal y5_re_DUT_out : std_logic_vector(31 downto 0);
  signal y5_im_DUT_out : std_logic_vector(31 downto 0);
  signal y6_re_DUT_out : std_logic_vector(31 downto 0);
  signal y6_im_DUT_out : std_logic_vector(31 downto 0);
  signal y7_re_DUT_out : std_logic_vector(31 downto 0);
  signal y7_im_DUT_out : std_logic_vector(31 downto 0);
  signal y8_re_DUT_out : std_logic_vector(31 downto 0);
  signal y8_im_DUT_out : std_logic_vector(31 downto 0);
  signal y9_re_DUT_out : std_logic_vector(31 downto 0);
  signal y9_im_DUT_out : std_logic_vector(31 downto 0);
  signal y10_re_DUT_out : std_logic_vector(31 downto 0);
  signal y10_im_DUT_out : std_logic_vector(31 downto 0);
  signal y11_re_DUT_out : std_logic_vector(31 downto 0);
  signal y11_im_DUT_out : std_logic_vector(31 downto 0);
  signal y12_re_DUT_out : std_logic_vector(31 downto 0);
  signal y12_im_DUT_out : std_logic_vector(31 downto 0);
  signal y13_re_DUT_out : std_logic_vector(31 downto 0);
  signal y13_im_DUT_out : std_logic_vector(31 downto 0);
  signal y14_re_DUT_out : std_logic_vector(31 downto 0);
  signal y14_im_DUT_out : std_logic_vector(31 downto 0);
  signal y15_re_DUT_out : std_logic_vector(31 downto 0);
  signal y15_im_DUT_out : std_logic_vector(31 downto 0);
  type output_mux_input_t is array (0 to 31) of std_logic_vector(31 downto 0);
  signal output_mux_input : output_mux_input_t;

  begin
    DUT : entity work.implementedSystem_toplevel
      port map (
        clk => clk,
        rst => rst,
        x0_re => x0_re_DUT_in,
        x0_im => x0_im_DUT_in,
        x1_re => x1_re_DUT_in,
        x1_im => x1_im_DUT_in,
        x2_re => x2_re_DUT_in,
        x2_im => x2_im_DUT_in,
        x3_re => x3_re_DUT_in,
        x3_im => x3_im_DUT_in,
        x4_re => x4_re_DUT_in,
        x4_im => x4_im_DUT_in,
        x5_re => x5_re_DUT_in,
        x5_im => x5_im_DUT_in,
        x6_re => x6_re_DUT_in,
        x6_im => x6_im_DUT_in,
        x7_re => x7_re_DUT_in,
        x7_im => x7_im_DUT_in,
        x8_re => x8_re_DUT_in,
        x8_im => x8_im_DUT_in,
        x9_re => x9_re_DUT_in,
        x9_im => x9_im_DUT_in,
        x10_re => x10_re_DUT_in,
        x10_im => x10_im_DUT_in,
        x11_re => x11_re_DUT_in,
        x11_im => x11_im_DUT_in,
        x12_re => x12_re_DUT_in,
        x12_im => x12_im_DUT_in,
        x13_re => x13_re_DUT_in,
        x13_im => x13_im_DUT_in,
        x14_re => x14_re_DUT_in,
        x14_im => x14_im_DUT_in,
        x15_re => x15_re_DUT_in,
        x15_im => x15_im_DUT_in,
        y0_re => y0_re_DUT_out,
        y0_im => y0_im_DUT_out,
        y1_re => y1_re_DUT_out,
        y1_im => y1_im_DUT_out,
        y2_re => y2_re_DUT_out,
        y2_im => y2_im_DUT_out,
        y3_re => y3_re_DUT_out,
        y3_im => y3_im_DUT_out,
        y4_re => y4_re_DUT_out,
        y4_im => y4_im_DUT_out,
        y5_re => y5_re_DUT_out,
        y5_im => y5_im_DUT_out,
        y6_re => y6_re_DUT_out,
        y6_im => y6_im_DUT_out,
        y7_re => y7_re_DUT_out,
        y7_im => y7_im_DUT_out,
        y8_re => y8_re_DUT_out,
        y8_im => y8_im_DUT_out,
        y9_re => y9_re_DUT_out,
        y9_im => y9_im_DUT_out,
        y10_re => y10_re_DUT_out,
        y10_im => y10_im_DUT_out,
        y11_re => y11_re_DUT_out,
        y11_im => y11_im_DUT_out,
        y12_re => y12_re_DUT_out,
        y12_im => y12_im_DUT_out,
        y13_re => y13_re_DUT_out,
        y13_im => y13_im_DUT_out,
        y14_re => y14_re_DUT_out,
        y14_im => y14_im_DUT_out,
        y15_re => y15_re_DUT_out,
        y15_im => y15_im_DUT_out
       );
    process(clk)
      begin
        if (rising_edge(clk)) then
          if (x0_re_enable = '1') then
            x0_re_DUT_in <= shared_input;
          end if; -- enable for input x0_re
          if (x0_im_enable = '1') then
            x0_im_DUT_in <= shared_input;
          end if; -- enable for input x0_im
          if (x1_re_enable = '1') then
            x1_re_DUT_in <= shared_input;
          end if; -- enable for input x1_re
          if (x1_im_enable = '1') then
            x1_im_DUT_in <= shared_input;
          end if; -- enable for input x1_im
          if (x2_re_enable = '1') then
            x2_re_DUT_in <= shared_input;
          end if; -- enable for input x2_re
          if (x2_im_enable = '1') then
            x2_im_DUT_in <= shared_input;
          end if; -- enable for input x2_im
          if (x3_re_enable = '1') then
            x3_re_DUT_in <= shared_input;
          end if; -- enable for input x3_re
          if (x3_im_enable = '1') then
            x3_im_DUT_in <= shared_input;
          end if; -- enable for input x3_im
          if (x4_re_enable = '1') then
            x4_re_DUT_in <= shared_input;
          end if; -- enable for input x4_re
          if (x4_im_enable = '1') then
            x4_im_DUT_in <= shared_input;
          end if; -- enable for input x4_im
          if (x5_re_enable = '1') then
            x5_re_DUT_in <= shared_input;
          end if; -- enable for input x5_re
          if (x5_im_enable = '1') then
            x5_im_DUT_in <= shared_input;
          end if; -- enable for input x5_im
          if (x6_re_enable = '1') then
            x6_re_DUT_in <= shared_input;
          end if; -- enable for input x6_re
          if (x6_im_enable = '1') then
            x6_im_DUT_in <= shared_input;
          end if; -- enable for input x6_im
          if (x7_re_enable = '1') then
            x7_re_DUT_in <= shared_input;
          end if; -- enable for input x7_re
          if (x7_im_enable = '1') then
            x7_im_DUT_in <= shared_input;
          end if; -- enable for input x7_im
          if (x8_re_enable = '1') then
            x8_re_DUT_in <= shared_input;
          end if; -- enable for input x8_re
          if (x8_im_enable = '1') then
            x8_im_DUT_in <= shared_input;
          end if; -- enable for input x8_im
          if (x9_re_enable = '1') then
            x9_re_DUT_in <= shared_input;
          end if; -- enable for input x9_re
          if (x9_im_enable = '1') then
            x9_im_DUT_in <= shared_input;
          end if; -- enable for input x9_im
          if (x10_re_enable = '1') then
            x10_re_DUT_in <= shared_input;
          end if; -- enable for input x10_re
          if (x10_im_enable = '1') then
            x10_im_DUT_in <= shared_input;
          end if; -- enable for input x10_im
          if (x11_re_enable = '1') then
            x11_re_DUT_in <= shared_input;
          end if; -- enable for input x11_re
          if (x11_im_enable = '1') then
            x11_im_DUT_in <= shared_input;
          end if; -- enable for input x11_im
          if (x12_re_enable = '1') then
            x12_re_DUT_in <= shared_input;
          end if; -- enable for input x12_re
          if (x12_im_enable = '1') then
            x12_im_DUT_in <= shared_input;
          end if; -- enable for input x12_im
          if (x13_re_enable = '1') then
            x13_re_DUT_in <= shared_input;
          end if; -- enable for input x13_re
          if (x13_im_enable = '1') then
            x13_im_DUT_in <= shared_input;
          end if; -- enable for input x13_im
          if (x14_re_enable = '1') then
            x14_re_DUT_in <= shared_input;
          end if; -- enable for input x14_re
          if (x14_im_enable = '1') then
            x14_im_DUT_in <= shared_input;
          end if; -- enable for input x14_im
          if (x15_re_enable = '1') then
            x15_re_DUT_in <= shared_input;
          end if; -- enable for input x15_re
          if (x15_im_enable = '1') then
            x15_im_DUT_in <= shared_input;
          end if; -- enable for input x15_im
        end if; -- clk
      end process;
    output_mux_input(0) <= y0_re_DUT_out;
    output_mux_input(1) <= y0_im_DUT_out;
    output_mux_input(2) <= y1_re_DUT_out;
    output_mux_input(3) <= y1_im_DUT_out;
    output_mux_input(4) <= y2_re_DUT_out;
    output_mux_input(5) <= y2_im_DUT_out;
    output_mux_input(6) <= y3_re_DUT_out;
    output_mux_input(7) <= y3_im_DUT_out;
    output_mux_input(8) <= y4_re_DUT_out;
    output_mux_input(9) <= y4_im_DUT_out;
    output_mux_input(10) <= y5_re_DUT_out;
    output_mux_input(11) <= y5_im_DUT_out;
    output_mux_input(12) <= y6_re_DUT_out;
    output_mux_input(13) <= y6_im_DUT_out;
    output_mux_input(14) <= y7_re_DUT_out;
    output_mux_input(15) <= y7_im_DUT_out;
    output_mux_input(16) <= y8_re_DUT_out;
    output_mux_input(17) <= y8_im_DUT_out;
    output_mux_input(18) <= y9_re_DUT_out;
    output_mux_input(19) <= y9_im_DUT_out;
    output_mux_input(20) <= y10_re_DUT_out;
    output_mux_input(21) <= y10_im_DUT_out;
    output_mux_input(22) <= y11_re_DUT_out;
    output_mux_input(23) <= y11_im_DUT_out;
    output_mux_input(24) <= y12_re_DUT_out;
    output_mux_input(25) <= y12_im_DUT_out;
    output_mux_input(26) <= y13_re_DUT_out;
    output_mux_input(27) <= y13_im_DUT_out;
    output_mux_input(28) <= y14_re_DUT_out;
    output_mux_input(29) <= y14_im_DUT_out;
    output_mux_input(30) <= y15_re_DUT_out;
    output_mux_input(31) <= y15_im_DUT_out;
    shared_output <= output_mux_input(to_integer(unsigned(output_select)));
    
end architecture;
