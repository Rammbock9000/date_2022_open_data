--------------------------------------------------------------------------------
--                         ModuloCounter_12_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity ModuloCounter_12_component is
   port ( clk, rst : in std_logic;
          Counter_out : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of ModuloCounter_12_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk,rst)
	 variable count : std_logic_vector(3 downto 0) := (others => '0');
begin
	 if rst = '1' then
	 	 count := (others => '0');
	 elsif clk'event and clk = '1' then
	 	 if count = 11 then
	 	 	 count := (others => '0');
	 	 else
	 	 	 count := count+1;
	 	 end if;
	 end if;
	 Counter_out <= count;
end process;
end architecture;

--------------------------------------------------------------------------------
--                          InputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2008)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity InputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(31 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of InputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal expInfty : std_logic := '0';
signal fracZero : std_logic := '0';
signal reprSubNormal : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal infinity : std_logic := '0';
signal zero : std_logic := '0';
signal NaN : std_logic := '0';
signal exnR : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   sX  <= X(31);
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   expInfty  <= '1' when expX = (7 downto 0 => '1') else '0';
   fracZero <= '1' when fracX = (22 downto 0 => '0') else '0';
   reprSubNormal <= fracX(22);
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= fracX(21 downto 0) & '0' when (expZero='1' and reprSubNormal='1')    else fracX;
   fracR <= sfracX;
   -- copy exponent. This will be OK even for subnormals, zero and infty since in such cases the exn bits will prevail
   expR <= expX;
   infinity <= expInfty and fracZero;
   zero <= expZero and not reprSubNormal;
   NaN <= expInfty and not fracZero;
   exnR <= 
           "00" when zero='1' 
      else "10" when infinity='1' 
      else "11" when NaN='1' 
      else "01" ;  -- normal number
   R <= exnR & sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--                         OutputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. Ferrandi  (2009-2012)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity OutputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of OutputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal exnX : std_logic_vector(1 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   exnX  <= X(33 downto 32);
   sX  <= X(31) when (exnX = "01" or exnX = "10" or exnX = "00") else '0';
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= 
      (22 downto 0 => '0') when (exnX = "00") else
      '1' & fracX(22 downto 1) when (expZero = '1' and exnX = "01") else
      fracX when (exnX = "01") else 
      (22 downto 1 => '0') & exnX(0);
   fracR <= sfracX;
   expR <=  
      (7 downto 0 => '0') when (exnX = "00") else
      expX when (exnX = "01") else 
      (7 downto 0 => '1');
   R <= sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_7_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_7_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(2 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_7_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000",
         iS_1 when "001",
         iS_2 when "010",
         iS_3 when "011",
         iS_4 when "100",
         iS_5 when "101",
         iS_6 when "110",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      Y <= s0;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid679703_RightShifter
--                 (RightShifter_24_by_max_26_F250_uid679705)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid679703_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid679703_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_27_f250_uid679708
--                  (IntAdderAlternative_27_f250_uid679712)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid679708 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid679708 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--               LZCShifter_28_to_28_counting_32_F250_uid679715
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid679715 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid679715 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_34_f250_uid679718
--                   (IntAdderClassical_34_f250_uid679720)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid679718 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid679718 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                            FPAdd_8_23_uid679703
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid679703 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid679703 is
   component FPAdd_8_23_uid679703_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid679708 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid679715 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid679718 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid679703_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid679708  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid679715  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid679718  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   component FPAdd_8_23_uid679703 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= Y;
   FPAddSubOp_instance: FPAdd_8_23_uid679703  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_12_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_12_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(3 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_12_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "0000",
         iS_1 when "0001",
         iS_2 when "0010",
         iS_3 when "0011",
         iS_4 when "0100",
         iS_5 when "0101",
         iS_6 when "0110",
         iS_7 when "0111",
         iS_8 when "1000",
         iS_9 when "1001",
         iS_10 when "1010",
         iS_11 when "1011",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_4_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(1 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "00",
         iS_1 when "01",
         iS_2 when "10",
         iS_3 when "11",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--          IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid681882
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid681882 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          Y : in std_logic_vector(23 downto 0);
          R : out std_logic_vector(47 downto 0)   );
end entity;

architecture arch of IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid681882 is
signal XX_m681883 : std_logic_vector(23 downto 0) := (others => '0');
signal YY_m681883 : std_logic_vector(23 downto 0) := (others => '0');
signal XX : unsigned(-1+24 downto 0) := (others => '0');
signal YY : unsigned(-1+24 downto 0) := (others => '0');
signal RR : unsigned(-1+48 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   XX_m681883 <= X ;
   YY_m681883 <= Y ;
   XX <= unsigned(X);
   YY <= unsigned(Y);
   RR <= XX*YY;
   R <= std_logic_vector(RR(47 downto 0));
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_33_f500_uid681886
--                   (IntAdderClassical_33_f500_uid681888)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_33_f500_uid681886 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(32 downto 0);
          Y : in std_logic_vector(32 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(32 downto 0)   );
end entity;

architecture arch of IntAdder_33_f500_uid681886 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--         FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin 2008-2011
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   component IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid681882 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             Y : in std_logic_vector(23 downto 0);
             R : out std_logic_vector(47 downto 0)   );
   end component;

   component IntAdder_33_f500_uid681886 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(32 downto 0);
             Y : in std_logic_vector(32 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(32 downto 0)   );
   end component;

signal sign, sign_d1, sign_d2 : std_logic := '0';
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal expY : std_logic_vector(7 downto 0) := (others => '0');
signal expSumPreSub, expSumPreSub_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal bias, bias_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal expSum : std_logic_vector(9 downto 0) := (others => '0');
signal sigX : std_logic_vector(23 downto 0) := (others => '0');
signal sigY : std_logic_vector(23 downto 0) := (others => '0');
signal sigProd, sigProd_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal excSel : std_logic_vector(3 downto 0) := (others => '0');
signal exc, exc_d1, exc_d2 : std_logic_vector(1 downto 0) := (others => '0');
signal norm : std_logic := '0';
signal expPostNorm : std_logic_vector(9 downto 0) := (others => '0');
signal sigProdExt, sigProdExt_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal expSig, expSig_d1 : std_logic_vector(32 downto 0) := (others => '0');
signal sticky, sticky_d1 : std_logic := '0';
signal guard, guard_d1 : std_logic := '0';
signal round : std_logic := '0';
signal expSigPostRound : std_logic_vector(32 downto 0) := (others => '0');
signal excPostNorm : std_logic_vector(1 downto 0) := (others => '0');
signal finalExc : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            sign_d1 <=  sign;
            sign_d2 <=  sign_d1;
            expSumPreSub_d1 <=  expSumPreSub;
            bias_d1 <=  bias;
            sigProd_d1 <=  sigProd;
            exc_d1 <=  exc;
            exc_d2 <=  exc_d1;
            sigProdExt_d1 <=  sigProdExt;
            expSig_d1 <=  expSig;
            sticky_d1 <=  sticky;
            guard_d1 <=  guard;
         end if;
      end process;
   sign <= X(31) xor Y(31);
   expX <= X(30 downto 23);
   expY <= Y(30 downto 23);
   expSumPreSub <= ("00" & expX) + ("00" & expY);
   bias <= CONV_STD_LOGIC_VECTOR(127,10);
   ----------------Synchro barrier, entering cycle 1----------------
   expSum <= expSumPreSub_d1 - bias_d1;
   ----------------Synchro barrier, entering cycle 0----------------
   sigX <= "1" & X(22 downto 0);
   sigY <= "1" & Y(22 downto 0);
   SignificandMultiplication: IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid681882  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => sigProd,
                 X => sigX,
                 Y => sigY);
   ----------------Synchro barrier, entering cycle 0----------------
   excSel <= X(33 downto 32) & Y(33 downto 32);
   with excSel select 
   exc <= "00" when  "0000" | "0001" | "0100", 
          "01" when "0101",
          "10" when "0110" | "1001" | "1010" ,
          "11" when others;
   norm <= sigProd_d1(47);
   -- exponent update
   expPostNorm <= expSum + ("000000000" & norm);
   -- significand normalization shift
   sigProdExt <= sigProd_d1(46 downto 0) & "0" when norm='1' else
                         sigProd_d1(45 downto 0) & "00";
   expSig <= expPostNorm & sigProdExt(47 downto 25);
   sticky <= sigProdExt(24);
   guard <= '0' when sigProdExt(23 downto 0)="000000000000000000000000" else '1';
   ----------------Synchro barrier, entering cycle 2----------------
   round <= sticky_d1 and ( (guard_d1 and not(sigProdExt_d1(25))) or (sigProdExt_d1(25) ))  ;
      RoundingAdder: IntAdder_33_f500_uid681886  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => round,
                 R => expSigPostRound,
                 X => expSig_d1,
                 Y => "000000000000000000000000000000000");
   with expSigPostRound(32 downto 31) select
   excPostNorm <=  "01"  when  "00",
                               "10"             when "01", 
                               "00"             when "11"|"10",
                               "11"             when others;
   with exc_d2 select 
   finalExc <= exc_d2 when  "11"|"10"|"00",
                       excPostNorm when others; 
   R <= finalExc & sign_d2 & expSigPostRound(30 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid682189_RightShifter
--                 (RightShifter_24_by_max_26_F250_uid682191)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid682189_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid682189_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_27_f250_uid682194
--                  (IntAdderAlternative_27_f250_uid682198)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid682194 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid682194 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--               LZCShifter_28_to_28_counting_32_F250_uid682201
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid682201 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid682201 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_34_f250_uid682204
--                   (IntAdderClassical_34_f250_uid682206)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid682204 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid682204 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                            FPAdd_8_23_uid682189
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid682189 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid682189 is
   component FPAdd_8_23_uid682189_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid682194 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid682201 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid682204 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid682189_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid682194  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid682201  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid682204  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
   component FPAdd_8_23_uid682189 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= (Y(Y'length-1 downto Y'length-2)) & (not Y(Y'length-3)) & Y(Y'length-4 downto 0);
   FPAddSubOp_instance: FPAdd_8_23_uid682189  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--                      Constant_float_8_23_1_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_1_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_1_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111100000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                      Constant_float_8_23_0_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_0_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_0_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0000000000000000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_cosnpi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosnpi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosnpi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_sinnpi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinnpi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinnpi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn3_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn3_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn3_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn3_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn3_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn3_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_cosnpi_div_2_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosnpi_div_2_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosnpi_div_2_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0000000000000000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_sinnpi_div_2_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinnpi_div_2_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinnpi_div_2_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111100000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn5_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn5_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn5_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn5_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn5_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn5_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn3_mult_pi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn3_mult_pi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn3_mult_pi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn3_mult_pi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn3_mult_pi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn3_mult_pi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn7_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn7_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn7_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn7_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn7_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn7_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_cosnpi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosnpi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosnpi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_sinnpi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinnpi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinnpi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      Y <= s1;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      Y <= s2;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "100" when "0000",
      "000" when "0001",
      "101" when "0010",
      "110" when "0011",
      "000" when "0100",
      "000" when "0101",
      "000" when "0110",
      "001" when "0111",
      "000" when "1000",
      "010" when "1001",
      "011" when "1010",
      "000" when "1011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "100" when "0000",
      "000" when "0001",
      "101" when "0010",
      "110" when "0011",
      "000" when "0100",
      "000" when "0101",
      "000" when "0110",
      "001" when "0111",
      "000" when "1000",
      "010" when "1001",
      "011" when "1010",
      "000" when "1011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "110" when "0000",
      "000" when "0001",
      "000" when "0010",
      "000" when "0011",
      "001" when "0100",
      "000" when "0101",
      "010" when "0110",
      "011" when "0111",
      "000" when "1000",
      "100" when "1001",
      "000" when "1010",
      "101" when "1011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "110" when "0000",
      "000" when "0001",
      "000" when "0010",
      "000" when "0011",
      "001" when "0100",
      "000" when "0101",
      "010" when "0110",
      "011" when "0111",
      "000" when "1000",
      "100" when "1001",
      "000" when "1010",
      "101" when "1011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "001" when "0001",
      "000" when "0010",
      "010" when "0011",
      "011" when "0100",
      "000" when "0101",
      "100" when "0110",
      "000" when "0111",
      "101" when "1000",
      "110" when "1001",
      "000" when "1010",
      "000" when "1011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "001" when "0001",
      "000" when "0010",
      "010" when "0011",
      "011" when "0100",
      "000" when "0101",
      "100" when "0110",
      "000" when "0111",
      "101" when "1000",
      "110" when "1001",
      "000" when "1010",
      "000" when "1011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "110" when "0000",
      "000" when "0001",
      "000" when "0010",
      "000" when "0011",
      "001" when "0100",
      "000" when "0101",
      "010" when "0110",
      "011" when "0111",
      "000" when "1000",
      "100" when "1001",
      "000" when "1010",
      "101" when "1011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "101" when "0000",
      "110" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "001" when "0101",
      "000" when "0110",
      "010" when "0111",
      "011" when "1000",
      "000" when "1001",
      "100" when "1010",
      "000" when "1011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "100" when "0000",
      "000" when "0001",
      "101" when "0010",
      "110" when "0011",
      "000" when "0100",
      "000" when "0101",
      "000" when "0110",
      "001" when "0111",
      "000" when "1000",
      "010" when "1001",
      "011" when "1010",
      "000" when "1011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "100" when "0000",
      "000" when "0001",
      "101" when "0010",
      "110" when "0011",
      "000" when "0100",
      "000" when "0101",
      "000" when "0110",
      "001" when "0111",
      "000" when "1000",
      "010" when "1001",
      "011" when "1010",
      "000" when "1011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "110" when "0000",
      "000" when "0001",
      "000" when "0010",
      "000" when "0011",
      "001" when "0100",
      "000" when "0101",
      "010" when "0110",
      "011" when "0111",
      "000" when "1000",
      "100" when "1001",
      "000" when "1010",
      "101" when "1011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "110" when "0000",
      "000" when "0001",
      "000" when "0010",
      "000" when "0011",
      "001" when "0100",
      "000" when "0101",
      "010" when "0110",
      "011" when "0111",
      "000" when "1000",
      "100" when "1001",
      "000" when "1010",
      "101" when "1011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "001" when "0001",
      "000" when "0010",
      "010" when "0011",
      "011" when "0100",
      "000" when "0101",
      "100" when "0110",
      "000" when "0111",
      "101" when "1000",
      "110" when "1001",
      "000" when "1010",
      "000" when "1011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "010" when "0001",
      "000" when "0010",
      "011" when "0011",
      "000" when "0100",
      "000" when "0101",
      "100" when "0110",
      "000" when "0111",
      "101" when "1000",
      "110" when "1001",
      "000" when "1010",
      "001" when "1011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "101" when "0000",
      "110" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "001" when "0101",
      "000" when "0110",
      "010" when "0111",
      "011" when "1000",
      "000" when "1001",
      "100" when "1010",
      "000" when "1011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "101" when "0000",
      "110" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "001" when "0101",
      "000" when "0110",
      "010" when "0111",
      "011" when "1000",
      "000" when "1001",
      "100" when "1010",
      "000" when "1011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "100" when "0000",
      "000" when "0001",
      "101" when "0010",
      "110" when "0011",
      "000" when "0100",
      "000" when "0101",
      "000" when "0110",
      "001" when "0111",
      "000" when "1000",
      "010" when "1001",
      "011" when "1010",
      "000" when "1011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "100" when "0000",
      "000" when "0001",
      "101" when "0010",
      "110" when "0011",
      "000" when "0100",
      "000" when "0101",
      "000" when "0110",
      "001" when "0111",
      "000" when "1000",
      "010" when "1001",
      "011" when "1010",
      "000" when "1011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "110" when "0000",
      "000" when "0001",
      "000" when "0010",
      "000" when "0011",
      "001" when "0100",
      "000" when "0101",
      "010" when "0110",
      "011" when "0111",
      "000" when "1000",
      "100" when "1001",
      "000" when "1010",
      "101" when "1011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "110" when "0000",
      "000" when "0001",
      "000" when "0010",
      "000" when "0011",
      "001" when "0100",
      "000" when "0101",
      "010" when "0110",
      "011" when "0111",
      "000" when "1000",
      "100" when "1001",
      "000" when "1010",
      "101" when "1011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "001" when "0001",
      "000" when "0010",
      "010" when "0011",
      "011" when "0100",
      "000" when "0101",
      "100" when "0110",
      "000" when "0111",
      "101" when "1000",
      "110" when "1001",
      "000" when "1010",
      "000" when "1011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "001" when "0001",
      "000" when "0010",
      "010" when "0011",
      "011" when "0100",
      "000" when "0101",
      "100" when "0110",
      "000" when "0111",
      "101" when "1000",
      "110" when "1001",
      "000" when "1010",
      "000" when "1011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "101" when "0000",
      "110" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "001" when "0101",
      "000" when "0110",
      "010" when "0111",
      "011" when "1000",
      "000" when "1001",
      "100" when "1010",
      "000" when "1011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "101" when "0000",
      "110" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "001" when "0101",
      "000" when "0110",
      "010" when "0111",
      "011" when "1000",
      "000" when "1001",
      "100" when "1010",
      "000" when "1011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "100" when "0000",
      "000" when "0001",
      "101" when "0010",
      "110" when "0011",
      "000" when "0100",
      "001" when "0101",
      "000" when "0110",
      "000" when "0111",
      "000" when "1000",
      "010" when "1001",
      "011" when "1010",
      "000" when "1011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "100" when "0000",
      "000" when "0001",
      "101" when "0010",
      "110" when "0011",
      "000" when "0100",
      "000" when "0101",
      "000" when "0110",
      "001" when "0111",
      "000" when "1000",
      "010" when "1001",
      "011" when "1010",
      "000" when "1011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "110" when "0000",
      "000" when "0001",
      "000" when "0010",
      "000" when "0011",
      "001" when "0100",
      "000" when "0101",
      "010" when "0110",
      "011" when "0111",
      "000" when "1000",
      "100" when "1001",
      "000" when "1010",
      "101" when "1011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "110" when "0000",
      "000" when "0001",
      "000" when "0010",
      "000" when "0011",
      "001" when "0100",
      "000" when "0101",
      "010" when "0110",
      "011" when "0111",
      "000" when "1000",
      "100" when "1001",
      "000" when "1010",
      "101" when "1011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "001" when "0001",
      "000" when "0010",
      "010" when "0011",
      "011" when "0100",
      "000" when "0101",
      "100" when "0110",
      "000" when "0111",
      "101" when "1000",
      "110" when "1001",
      "000" when "1010",
      "000" when "1011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "001" when "0001",
      "000" when "0010",
      "010" when "0011",
      "011" when "0100",
      "000" when "0101",
      "100" when "0110",
      "000" when "0111",
      "101" when "1000",
      "110" when "1001",
      "000" when "1010",
      "000" when "1011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "110" when "0001",
      "000" when "0010",
      "010" when "0011",
      "000" when "0100",
      "011" when "0101",
      "000" when "0110",
      "100" when "0111",
      "101" when "1000",
      "000" when "1001",
      "001" when "1010",
      "000" when "1011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "101" when "0000",
      "110" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "001" when "0101",
      "000" when "0110",
      "010" when "0111",
      "011" when "1000",
      "000" when "1001",
      "100" when "1010",
      "000" when "1011",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Add130_6_impl_0_LUT_wIn_4_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add130_6_impl_0_LUT_wIn_4_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add130_6_impl_0_LUT_wIn_4_wOut_2 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "00" when "0000",
      "11" when "0001",
      "00" when "0010",
      "00" when "0011",
      "00" when "0100",
      "00" when "0101",
      "10" when "0110",
      "00" when "0111",
      "01" when "1000",
      "00" when "1001",
      "00" when "1010",
      "00" when "1011",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Add130_6_impl_0_LUT_wIn_4_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add130_6_impl_0_LUT_wIn_4_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add130_6_impl_0_LUT_wIn_4_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Add130_6_impl_0_LUT_wIn_4_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Add130_6_impl_0_LUT_wIn_4_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Add130_6_impl_1_LUT_wIn_4_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add130_6_impl_1_LUT_wIn_4_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add130_6_impl_1_LUT_wIn_4_wOut_2 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "00" when "0000",
      "11" when "0001",
      "00" when "0010",
      "00" when "0011",
      "00" when "0100",
      "00" when "0101",
      "10" when "0110",
      "00" when "0111",
      "01" when "1000",
      "00" when "1001",
      "00" when "1010",
      "00" when "1011",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Add130_6_impl_1_LUT_wIn_4_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add130_6_impl_1_LUT_wIn_4_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add130_6_impl_1_LUT_wIn_4_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Add130_6_impl_1_LUT_wIn_4_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Add130_6_impl_1_LUT_wIn_4_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--        GenericLut_LUTData_MUX_Subtract125_6_impl_0_LUT_wIn_4_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract125_6_impl_0_LUT_wIn_4_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract125_6_impl_0_LUT_wIn_4_wOut_2 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "00" when "0000",
      "10" when "0001",
      "00" when "0010",
      "00" when "0011",
      "00" when "0100",
      "00" when "0101",
      "01" when "0110",
      "00" when "0111",
      "11" when "1000",
      "00" when "1001",
      "00" when "1010",
      "00" when "1011",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Subtract125_6_impl_0_LUT_wIn_4_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract125_6_impl_0_LUT_wIn_4_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract125_6_impl_0_LUT_wIn_4_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Subtract125_6_impl_0_LUT_wIn_4_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Subtract125_6_impl_0_LUT_wIn_4_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--        GenericLut_LUTData_MUX_Subtract125_6_impl_1_LUT_wIn_4_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract125_6_impl_1_LUT_wIn_4_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract125_6_impl_1_LUT_wIn_4_wOut_2 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "00" when "0000",
      "01" when "0001",
      "00" when "0010",
      "00" when "0011",
      "00" when "0100",
      "00" when "0101",
      "10" when "0110",
      "00" when "0111",
      "11" when "1000",
      "00" when "1001",
      "00" when "1010",
      "00" when "1011",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Subtract125_6_impl_1_LUT_wIn_4_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract125_6_impl_1_LUT_wIn_4_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract125_6_impl_1_LUT_wIn_4_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Subtract125_6_impl_1_LUT_wIn_4_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Subtract125_6_impl_1_LUT_wIn_4_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      Y <= s3;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 14 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      Y <= s13;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      Y <= s5;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 7 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      Y <= s6;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 9 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      Y <= s8;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 5 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      Y <= s4;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 15 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      Y <= s14;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 8 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      Y <= s7;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      Y <= s10;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 10 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      Y <= s9;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 20 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      Y <= s19;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 16 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      Y <= s15;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 13 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      Y <= s12;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 17 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      Y <= s16;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                         implementedSystem_toplevel
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity implementedSystem_toplevel is
   port ( clk, rst : in std_logic;
          x0_re_0 : in std_logic_vector(31 downto 0);
          x0_im_0 : in std_logic_vector(31 downto 0);
          x1_re_0 : in std_logic_vector(31 downto 0);
          x1_im_0 : in std_logic_vector(31 downto 0);
          x2_re_0 : in std_logic_vector(31 downto 0);
          x2_im_0 : in std_logic_vector(31 downto 0);
          x3_re_0 : in std_logic_vector(31 downto 0);
          x3_im_0 : in std_logic_vector(31 downto 0);
          x4_re_0 : in std_logic_vector(31 downto 0);
          x4_im_0 : in std_logic_vector(31 downto 0);
          x5_re_0 : in std_logic_vector(31 downto 0);
          x5_im_0 : in std_logic_vector(31 downto 0);
          x6_re_0 : in std_logic_vector(31 downto 0);
          x6_im_0 : in std_logic_vector(31 downto 0);
          x7_re_0 : in std_logic_vector(31 downto 0);
          x7_im_0 : in std_logic_vector(31 downto 0);
          x8_re_0 : in std_logic_vector(31 downto 0);
          x8_im_0 : in std_logic_vector(31 downto 0);
          x9_re_0 : in std_logic_vector(31 downto 0);
          x9_im_0 : in std_logic_vector(31 downto 0);
          x10_re_0 : in std_logic_vector(31 downto 0);
          x10_im_0 : in std_logic_vector(31 downto 0);
          x11_re_0 : in std_logic_vector(31 downto 0);
          x11_im_0 : in std_logic_vector(31 downto 0);
          x12_re_0 : in std_logic_vector(31 downto 0);
          x12_im_0 : in std_logic_vector(31 downto 0);
          x13_re_0 : in std_logic_vector(31 downto 0);
          x13_im_0 : in std_logic_vector(31 downto 0);
          x14_re_0 : in std_logic_vector(31 downto 0);
          x14_im_0 : in std_logic_vector(31 downto 0);
          x15_re_0 : in std_logic_vector(31 downto 0);
          x15_im_0 : in std_logic_vector(31 downto 0);
          y0_re_0 : out std_logic_vector(31 downto 0);
          y0_im_0 : out std_logic_vector(31 downto 0);
          y1_re_0 : out std_logic_vector(31 downto 0);
          y1_im_0 : out std_logic_vector(31 downto 0);
          y2_re_0 : out std_logic_vector(31 downto 0);
          y2_im_0 : out std_logic_vector(31 downto 0);
          y3_re_0 : out std_logic_vector(31 downto 0);
          y3_im_0 : out std_logic_vector(31 downto 0);
          y4_re_0 : out std_logic_vector(31 downto 0);
          y4_im_0 : out std_logic_vector(31 downto 0);
          y5_re_0 : out std_logic_vector(31 downto 0);
          y5_im_0 : out std_logic_vector(31 downto 0);
          y6_re_0 : out std_logic_vector(31 downto 0);
          y6_im_0 : out std_logic_vector(31 downto 0);
          y7_re_0 : out std_logic_vector(31 downto 0);
          y7_im_0 : out std_logic_vector(31 downto 0);
          y8_re_0 : out std_logic_vector(31 downto 0);
          y8_im_0 : out std_logic_vector(31 downto 0);
          y9_re_0 : out std_logic_vector(31 downto 0);
          y9_im_0 : out std_logic_vector(31 downto 0);
          y10_re_0 : out std_logic_vector(31 downto 0);
          y10_im_0 : out std_logic_vector(31 downto 0);
          y11_re_0 : out std_logic_vector(31 downto 0);
          y11_im_0 : out std_logic_vector(31 downto 0);
          y12_re_0 : out std_logic_vector(31 downto 0);
          y12_im_0 : out std_logic_vector(31 downto 0);
          y13_re_0 : out std_logic_vector(31 downto 0);
          y13_im_0 : out std_logic_vector(31 downto 0);
          y14_re_0 : out std_logic_vector(31 downto 0);
          y14_im_0 : out std_logic_vector(31 downto 0);
          y15_re_0 : out std_logic_vector(31 downto 0);
          y15_im_0 : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of implementedSystem_toplevel is
   component ModuloCounter_12_component is
      port ( clk, rst : in std_logic;
             Counter_out : out std_logic_vector(3 downto 0)   );
   end component;

   component InputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(31 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component OutputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(31 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_7_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(2 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_12_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(3 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_4_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(1 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_1_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_0_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosnpi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinnpi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn3_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn3_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosnpi_div_2_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinnpi_div_2_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn5_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn5_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn3_mult_pi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn3_mult_pi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn7_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn7_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosnpi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinnpi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add130_6_impl_0_LUT_wIn_4_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add130_6_impl_1_LUT_wIn_4_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Subtract125_6_impl_0_LUT_wIn_4_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Subtract125_6_impl_1_LUT_wIn_4_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

signal ModCount121_out : std_logic_vector(3 downto 0) := (others => '0');
signal x0_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x0_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x1_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x1_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x2_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x2_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x3_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x3_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x4_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x4_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x5_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x5_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x6_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x6_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x7_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x7_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x8_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x8_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x9_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x9_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x10_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x10_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x11_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x11_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x12_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x12_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x13_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x13_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x14_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x14_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x15_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x15_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y0_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y0_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y1_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y1_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y2_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y2_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y3_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y3_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y4_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y4_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y5_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y5_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y6_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y6_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y7_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No14_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y7_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No15_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y8_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No16_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y8_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No17_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y9_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No18_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y9_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No19_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y10_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No20_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y10_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No21_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y11_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No22_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y11_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No23_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y12_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No24_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y12_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No25_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y13_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No26_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y13_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No27_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y14_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No28_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y14_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No29_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y15_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No30_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y15_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No31_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No32_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No33_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No34_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No35_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No36_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No37_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No38_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No39_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No40_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No41_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No42_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No43_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No44_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No45_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No46_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No47_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No48_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No49_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No50_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No51_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No52_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No53_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No54_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No55_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No56_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No57_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No58_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No59_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add3_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No60_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No61_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add3_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No62_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No63_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add3_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No64_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No65_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add3_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No66_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No67_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add3_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No68_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No69_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add3_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No70_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No71_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add3_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No72_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No73_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add12_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No74_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No75_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add12_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No76_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No77_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add12_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No78_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No79_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add12_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No80_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No81_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add12_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No82_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No83_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add12_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No84_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No85_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add12_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No86_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No87_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add5_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add5_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No88_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add5_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No89_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add5_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add5_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No90_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add5_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No91_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add5_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add5_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No92_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add5_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No93_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add5_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add5_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No94_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add5_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No95_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add14_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add14_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No96_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add14_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No97_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add14_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add14_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No98_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add14_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No99_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add6_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add6_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No100_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add6_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No101_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add15_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add15_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No102_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add15_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No103_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add8_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add8_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No104_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add8_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No105_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add8_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add8_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No106_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add8_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No107_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add8_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add8_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No108_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add8_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No109_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add8_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add8_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No110_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add8_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No111_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add10_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add10_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No112_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add10_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No113_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add23_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add23_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No114_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add23_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No115_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add23_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add23_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No116_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add23_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No117_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add23_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add23_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No118_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add23_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No119_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add113_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add113_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No120_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add113_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No121_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add113_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add113_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No122_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add113_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No123_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add113_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add113_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No124_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add113_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No125_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add113_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add113_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No126_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add113_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No127_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add113_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add113_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No128_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add113_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No129_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add24_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add24_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No130_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add24_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No131_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add32_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add32_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No132_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add32_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No133_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add122_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add122_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No134_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add122_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No135_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add33_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add33_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No136_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add33_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No137_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add33_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add33_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No138_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add33_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No139_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add33_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add33_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No140_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add33_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No141_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add33_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add33_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No142_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add33_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No143_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add33_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add33_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No144_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add33_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No145_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add123_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add123_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No146_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add123_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No147_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add123_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add123_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No148_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add123_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No149_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add123_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add123_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No150_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add123_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No151_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add123_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add123_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No152_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add123_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No153_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add123_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add123_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No154_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add123_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No155_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add35_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add35_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No156_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add35_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No157_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add35_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add35_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No158_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add35_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No159_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add35_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add35_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No160_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add35_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No161_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add130_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add130_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No162_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add130_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No163_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No164_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No165_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No166_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No167_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No168_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No169_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No170_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No171_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No172_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No173_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No174_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No175_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No176_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No177_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No178_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No179_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No180_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No181_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No182_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No183_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No184_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No185_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No186_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No187_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No188_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No189_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No190_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No191_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No192_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No193_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No194_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No195_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No196_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No197_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No198_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No199_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No200_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No201_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No202_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No203_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No204_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No205_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product5_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product5_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No206_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product5_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No207_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product5_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product5_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No208_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product5_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No209_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product5_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product5_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No210_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product5_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No211_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product5_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product5_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No212_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product5_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No213_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product5_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product5_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No214_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product5_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No215_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product5_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product5_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No216_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product5_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No217_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product5_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product5_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No218_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product5_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No219_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product12_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No220_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No221_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product12_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No222_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No223_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product12_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No224_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No225_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product12_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No226_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No227_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product12_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No228_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No229_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product12_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No230_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No231_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product12_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No232_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No233_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product22_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product22_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No234_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product22_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No235_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product22_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product22_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No236_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product22_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No237_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product22_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product22_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No238_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product22_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No239_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product22_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product22_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No240_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product22_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No241_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product22_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product22_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No242_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product22_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No243_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product22_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product22_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No244_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product22_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No245_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product22_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product22_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No246_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product22_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No247_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No248_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No249_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No250_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No251_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No252_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No253_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No254_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No255_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No256_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No257_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No258_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No259_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No260_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No261_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract3_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No262_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No263_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract3_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No264_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No265_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract3_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No266_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No267_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract3_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No268_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No269_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract3_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No270_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No271_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract3_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No272_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No273_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract3_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No274_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No275_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product6_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No276_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No277_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product6_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No278_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No279_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product6_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No280_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No281_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product6_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No282_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No283_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product6_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No284_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No285_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product6_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No286_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No287_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product6_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No288_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No289_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product23_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No290_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No291_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product23_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No292_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No293_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product23_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No294_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No295_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product23_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No296_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No297_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product23_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No298_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No299_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product23_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No300_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No301_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product23_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No302_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No303_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product33_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No304_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No305_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product33_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No306_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No307_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product33_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No308_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No309_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product33_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No310_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No311_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product33_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No312_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No313_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product33_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No314_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No315_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product33_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No316_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No317_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract4_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No318_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No319_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract4_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No320_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No321_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract4_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No322_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No323_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract4_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No324_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No325_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract4_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No326_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No327_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract4_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No328_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No329_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract4_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No330_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No331_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract5_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract5_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No332_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract5_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No333_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract5_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract5_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No334_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract5_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No335_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product26_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product26_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No336_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product26_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No337_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product26_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product26_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No338_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product26_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No339_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product26_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product26_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No340_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product26_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No341_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product26_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product26_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No342_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product26_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No343_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product26_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product26_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No344_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product26_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No345_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product26_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product26_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No346_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product26_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No347_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product26_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product26_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No348_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product26_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No349_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract7_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract7_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No350_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract7_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No351_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract7_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract7_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No352_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract7_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No353_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract7_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract7_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No354_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract7_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No355_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract7_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract7_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No356_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract7_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No357_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract7_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract7_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No358_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract7_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No359_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract8_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract8_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No360_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract8_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No361_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract8_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract8_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No362_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract8_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No363_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract8_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract8_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No364_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract8_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No365_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract8_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract8_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No366_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract8_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No367_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product18_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product18_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No368_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product18_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No369_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product18_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product18_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No370_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product18_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No371_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product18_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product18_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No372_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product18_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No373_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product18_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product18_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No374_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product18_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No375_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product18_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product18_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No376_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product18_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No377_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product18_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product18_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No378_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product18_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No379_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product18_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product18_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No380_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product18_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No381_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product28_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No382_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No383_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product28_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No384_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No385_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product28_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No386_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No387_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product28_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No388_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No389_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product28_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No390_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No391_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product28_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No392_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No393_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product28_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No394_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No395_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract9_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No396_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No397_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract9_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No398_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No399_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract9_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No400_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No401_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract9_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No402_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No403_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract9_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No404_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No405_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract9_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No406_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No407_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract9_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No408_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No409_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract10_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract10_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No410_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract10_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No411_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product50_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product50_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No412_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product50_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No413_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product50_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product50_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No414_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product50_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No415_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product50_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product50_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No416_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product50_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No417_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product50_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product50_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No418_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product50_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No419_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product50_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product50_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No420_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product50_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No421_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product50_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product50_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No422_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product50_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No423_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product50_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product50_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No424_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product50_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No425_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product122_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product122_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No426_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product122_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No427_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product122_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product122_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No428_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product122_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No429_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product122_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product122_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No430_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product122_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No431_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product122_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product122_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No432_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product122_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No433_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product122_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product122_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No434_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product122_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No435_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product122_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product122_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No436_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product122_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No437_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product122_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product122_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No438_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product122_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No439_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product221_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product221_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No440_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product221_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No441_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product221_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product221_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No442_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product221_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No443_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product221_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product221_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No444_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product221_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No445_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product221_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product221_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No446_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product221_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No447_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product221_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product221_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No448_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product221_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No449_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product221_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product221_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No450_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product221_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No451_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product221_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product221_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No452_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product221_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No453_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product321_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No454_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No455_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product321_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No456_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No457_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product321_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No458_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No459_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product321_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No460_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No461_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product321_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No462_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No463_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product321_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No464_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No465_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product321_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No466_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No467_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract23_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract23_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No468_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract23_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No469_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract23_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract23_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No470_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract23_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No471_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract23_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract23_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No472_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract23_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No473_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract23_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract23_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No474_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract23_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No475_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract23_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract23_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No476_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract23_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No477_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract23_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract23_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No478_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract23_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No479_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract23_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract23_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No480_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract23_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No481_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract30_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract30_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No482_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract30_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No483_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract30_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract30_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No484_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract30_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No485_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract30_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract30_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No486_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract30_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No487_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract30_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract30_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No488_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract30_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No489_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract30_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract30_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No490_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract30_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No491_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract30_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract30_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No492_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract30_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No493_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract30_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract30_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No494_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract30_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No495_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract32_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract32_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No496_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract32_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No497_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract32_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract32_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No498_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract32_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No499_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract32_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract32_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No500_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract32_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No501_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract32_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract32_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No502_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract32_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No503_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract32_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract32_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No504_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract32_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No505_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract32_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract32_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No506_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract32_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No507_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract43_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract43_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No508_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract43_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No509_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract44_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract44_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No510_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract44_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No511_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract49_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract49_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No512_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract49_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No513_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract116_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract116_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No514_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract116_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No515_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract58_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract58_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No516_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract58_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No517_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract125_6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract125_6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No518_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract125_6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No519_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant2_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant11_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant4_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant13_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant5_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant14_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant6_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant15_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant7_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant16_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant8_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant17_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant9_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant18_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant1_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No168_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No169_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No170_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No171_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No172_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No173_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No174_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No182_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No183_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No184_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No185_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No186_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No187_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No188_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No210_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No211_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No212_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No213_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No214_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No215_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No216_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No217_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No218_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No219_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No220_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No221_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No222_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No223_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No224_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No225_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No226_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No227_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No228_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No229_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No230_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No238_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No239_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No240_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No241_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No242_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No243_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No244_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No259_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No260_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No261_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No262_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No263_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No264_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No265_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No266_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No267_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No268_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No269_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No270_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No271_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No272_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No14_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No15_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No16_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No17_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No18_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No19_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No20_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No42_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No43_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No44_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No45_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No46_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No47_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No48_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No42_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No43_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No44_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No45_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No46_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No47_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No48_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y0_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y0_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y1_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y1_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y2_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y2_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y3_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y3_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y4_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y4_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y5_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y5_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y6_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y6_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y7_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y7_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y8_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y8_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y9_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y9_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y10_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y10_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y11_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y11_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y12_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y12_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y13_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y13_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y14_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y14_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y15_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y15_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Add130_6_impl_0_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Add130_6_impl_1_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Subtract125_6_impl_0_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Subtract125_6_impl_1_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal SharedReg_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg360_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg408_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg434_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg463_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg465_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg470_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg477_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg481_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg483_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg485_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg500_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg508_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg510_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg512_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg528_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg531_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg533_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg534_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg536_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg582_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg587_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg588_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg592_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg601_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg602_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg604_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg605_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg607_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg616_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg620_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg626_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg629_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg634_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg644_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg646_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg649_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg666_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg667_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg670_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg676_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg680_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg681_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg682_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg688_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg690_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg702_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg703_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg705_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg706_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg721_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg724_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg725_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg731_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg736_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg740_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg745_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg750_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg751_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg756_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg757_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg761_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg762_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg763_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg765_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg771_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg774_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg775_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg823_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg844_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg864_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg869_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg870_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg873_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg874_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg875_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg877_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg878_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg879_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg880_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg881_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg890_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg891_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg892_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg893_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg894_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg895_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg896_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg897_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg898_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg905_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg915_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg919_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg923_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg925_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg930_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg944_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg945_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg946_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg949_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg950_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg951_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg952_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg953_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg954_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg955_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg956_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg958_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg959_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg960_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg961_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg962_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg963_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg964_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg965_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg966_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg967_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg969_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg970_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg971_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg972_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg973_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg974_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg975_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg976_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg977_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg978_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg979_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg980_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg981_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg982_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg983_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg984_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg985_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg986_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg987_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg988_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg989_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg990_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg991_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg992_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg993_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg994_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg995_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg996_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg997_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg999_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1000_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1001_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1002_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1003_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1004_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1005_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1006_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1007_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1008_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1009_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1010_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1012_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1013_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1014_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1015_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1016_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1017_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1018_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1019_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1020_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1021_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1022_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1023_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1024_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1025_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1026_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1028_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1029_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1030_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1031_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1032_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1033_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1034_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1035_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1036_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1038_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1039_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1040_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1041_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1042_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1043_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1044_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1045_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1046_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1047_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1048_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1049_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1050_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1051_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1052_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1053_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1054_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1055_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1056_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1058_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1059_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1060_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1061_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1062_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1064_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1065_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1066_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1067_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1068_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1069_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1070_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1071_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1072_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1073_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1074_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1075_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1077_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1078_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1079_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1080_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1081_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1082_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1083_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1084_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1085_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1087_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1088_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1089_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1090_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1091_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1092_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1093_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1094_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1095_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1096_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1097_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1098_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1099_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1100_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1101_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1102_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1105_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1127_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1128_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1130_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1132_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1133_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1138_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1142_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1143_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1144_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1145_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1146_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1147_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1148_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1149_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1150_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1151_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1153_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1154_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1155_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1156_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1157_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1159_out : std_logic_vector(33 downto 0) := (others => '0');
signal x0_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x0_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x1_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x1_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x2_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x2_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x3_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x3_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x4_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x4_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x5_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x5_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x6_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x6_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x7_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x7_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x8_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x8_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x9_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x9_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x10_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x10_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x11_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x11_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x12_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x12_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x13_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x13_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x14_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x14_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x15_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x15_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y0_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y0_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y1_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y1_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y2_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y2_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y3_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y3_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y4_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y4_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y5_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y5_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y6_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y6_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y7_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y7_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y8_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1042_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1047_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1054_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1022_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1028_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1066_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y8_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg1070_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1081_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1060_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1075_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y9_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg1004_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg984_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg986_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg990_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg993_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1028_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1033_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y9_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1007_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1012_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1017_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1022_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1060_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1066_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y10_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg666_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y10_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y11_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg1004_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg984_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg986_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1017_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg993_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg997_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1066_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y11_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1007_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1012_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1054_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1022_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1028_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1075_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y12_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1094_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1088_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y12_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg981_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg984_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg986_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg990_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1001_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y13_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg1070_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1042_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1047_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1054_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1075_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y13_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg1094_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1081_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1088_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y14_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg981_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1001_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y14_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg1004_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg984_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg997_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1033_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y15_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg1060_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1070_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1042_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1047_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1088_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y15_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg1094_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1081_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1101_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No32_out_to_Add2_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No33_out_to_Add2_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1004_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg666_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg982_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No34_out_to_Add2_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No35_out_to_Add2_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No1_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1009_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1084_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1007_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No36_out_to_Add2_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No37_out_to_Add2_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1014_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg879_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg986_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No38_out_to_Add2_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No39_out_to_Add2_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg877_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No3_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1017_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No3_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No40_out_to_Add2_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No41_out_to_Add2_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg705_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1023_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg705_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No4_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No42_out_to_Add2_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No43_out_to_Add2_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg997_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg930_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg952_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg996_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No263_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No44_out_to_Add2_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No45_out_to_Add2_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg874_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1033_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg360_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg997_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg976_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No6_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1032_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1002_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg954_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No46_out_to_Add11_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No47_out_to_Add11_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1006_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1073_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg434_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg667_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No48_out_to_Add11_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No49_out_to_Add11_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg676_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg483_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No50_out_to_Add11_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No51_out_to_Add11_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No2_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No2_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No52_out_to_Add11_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No53_out_to_Add11_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1055_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No54_out_to_Add11_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No55_out_to_Add11_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg587_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg706_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg763_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No56_out_to_Add11_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No57_out_to_Add11_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg470_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg973_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg765_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No5_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg951_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No58_out_to_Add11_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No59_out_to_Add11_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1035_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1078_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg771_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg703_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg602_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No60_out_to_Add3_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No61_out_to_Add3_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg481_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No62_out_to_Add3_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No63_out_to_Add3_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1044_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No64_out_to_Add3_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No65_out_to_Add3_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg682_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1049_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No66_out_to_Add3_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No67_out_to_Add3_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg582_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg991_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No68_out_to_Add3_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No69_out_to_Add3_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No4_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg994_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg463_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No70_out_to_Add3_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No71_out_to_Add3_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1030_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg592_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg869_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No72_out_to_Add3_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No73_out_to_Add3_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1066_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No74_out_to_Add12_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No75_out_to_Add12_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1039_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg481_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg670_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No76_out_to_Add12_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No77_out_to_Add12_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No1_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg985_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg775_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No78_out_to_Add12_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No79_out_to_Add12_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg681_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No2_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg987_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No80_out_to_Add12_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No81_out_to_Add12_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg864_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No3_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg923_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg881_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No82_out_to_Add12_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No83_out_to_Add12_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg588_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg616_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg951_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No84_out_to_Add12_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No85_out_to_Add12_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No5_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No86_out_to_Add12_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No87_out_to_Add12_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1068_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg873_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg875_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No88_out_to_Add5_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No89_out_to_Add5_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg962_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1007_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No90_out_to_Add5_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No91_out_to_Add5_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg964_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg965_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg750_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1012_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No260_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No92_out_to_Add5_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No93_out_to_Add5_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Add5_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg986_out_to_MUX_Add5_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Add5_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg919_out_to_MUX_Add5_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No219_out_to_MUX_Add5_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add5_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out_to_MUX_Add5_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Add5_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Add5_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg880_out_to_MUX_Add5_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1017_out_to_MUX_Add5_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Add5_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Add5_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg989_out_to_MUX_Add5_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Add5_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg892_out_to_MUX_Add5_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No226_out_to_MUX_Add5_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add5_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Add5_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out_to_MUX_Add5_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg946_out_to_MUX_Add5_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out_to_MUX_Add5_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_Add5_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Add5_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No94_out_to_Add5_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No95_out_to_Add5_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Add5_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Add5_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg705_out_to_MUX_Add5_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out_to_MUX_Add5_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg970_out_to_MUX_Add5_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out_to_MUX_Add5_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add5_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg731_out_to_MUX_Add5_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg971_out_to_MUX_Add5_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add5_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Add5_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out_to_MUX_Add5_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Add5_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Add5_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out_to_MUX_Add5_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Add5_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Add5_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No262_out_to_MUX_Add5_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add5_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out_to_MUX_Add5_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out_to_MUX_Add5_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add5_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Add5_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out_to_MUX_Add5_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No96_out_to_Add14_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No97_out_to_Add14_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Add14_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out_to_MUX_Add14_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Add14_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1061_out_to_MUX_Add14_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Add14_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Add14_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Add14_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Add14_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out_to_MUX_Add14_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out_to_MUX_Add14_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add14_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add14_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out_to_MUX_Add14_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Add14_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_Add14_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_Add14_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Add14_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Add14_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Add14_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Add14_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out_to_MUX_Add14_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Add14_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add14_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add14_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No98_out_to_Add14_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No99_out_to_Add14_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Add14_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No6_out_to_MUX_Add14_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Add14_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg703_out_to_MUX_Add14_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Add14_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out_to_MUX_Add14_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Add14_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out_to_MUX_Add14_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Add14_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg745_out_to_MUX_Add14_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Add14_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add14_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add14_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Add14_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_Add14_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1002_out_to_MUX_Add14_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Add14_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Add14_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Add14_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Add14_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Add14_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No188_out_to_MUX_Add14_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out_to_MUX_Add14_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add14_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No100_out_to_Add6_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No101_out_to_Add6_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg993_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg990_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg923_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No220_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No45_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg761_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg949_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg992_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg896_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No227_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg634_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg925_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg949_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No102_out_to_Add15_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No103_out_to_Add15_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Add15_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Add15_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Add15_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg967_out_to_MUX_Add15_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out_to_MUX_Add15_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add15_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Add15_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add15_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out_to_MUX_Add15_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg688_out_to_MUX_Add15_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Add15_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1019_out_to_MUX_Add15_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Add15_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Add15_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Add15_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg945_out_to_MUX_Add15_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No261_out_to_MUX_Add15_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add15_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Add15_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add15_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out_to_MUX_Add15_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Add15_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Add15_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg757_out_to_MUX_Add15_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No104_out_to_Add8_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No105_out_to_Add8_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out_to_MUX_Add8_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add8_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add8_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No_out_to_MUX_Add8_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out_to_MUX_Add8_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out_to_MUX_Add8_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Add8_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Add8_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Add8_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg981_out_to_MUX_Add8_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Add8_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg721_out_to_MUX_Add8_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out_to_MUX_Add8_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add8_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add8_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Add8_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Add8_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg982_out_to_MUX_Add8_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Add8_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg666_out_to_MUX_Add8_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Add8_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_Add8_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Add8_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No182_out_to_MUX_Add8_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No106_out_to_Add8_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No107_out_to_Add8_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Add8_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out_to_MUX_Add8_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Add8_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out_to_MUX_Add8_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out_to_MUX_Add8_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Add8_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Add8_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Add8_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add8_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Add8_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out_to_MUX_Add8_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Add8_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out_to_MUX_Add8_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Add8_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_Add8_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_Add8_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg762_out_to_MUX_Add8_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Add8_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Add8_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Add8_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add8_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add8_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Add8_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg616_out_to_MUX_Add8_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No108_out_to_Add8_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No109_out_to_Add8_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Add8_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Add8_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Add8_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Add8_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out_to_MUX_Add8_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Add8_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Add8_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Add8_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Add8_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out_to_MUX_Add8_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add8_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Add8_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Add8_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg954_out_to_MUX_Add8_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out_to_MUX_Add8_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Add8_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out_to_MUX_Add8_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_Add8_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Add8_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Add8_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Add8_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Add8_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add8_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add8_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No110_out_to_Add8_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No111_out_to_Add8_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Add8_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Add8_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Add8_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out_to_MUX_Add8_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out_to_MUX_Add8_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Add8_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg702_out_to_MUX_Add8_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Add8_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Add8_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No244_out_to_MUX_Add8_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out_to_MUX_Add8_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add8_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg745_out_to_MUX_Add8_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out_to_MUX_Add8_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out_to_MUX_Add8_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out_to_MUX_Add8_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out_to_MUX_Add8_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Add8_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Add8_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Add8_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out_to_MUX_Add8_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Add8_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Add8_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add8_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No112_out_to_Add10_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No113_out_to_Add10_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add10_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Add10_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg477_out_to_MUX_Add10_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Add10_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out_to_MUX_Add10_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Add10_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Add10_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out_to_MUX_Add10_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Add10_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Add10_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add10_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Add10_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add10_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg955_out_to_MUX_Add10_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out_to_MUX_Add10_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg954_out_to_MUX_Add10_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Add10_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg955_out_to_MUX_Add10_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Add10_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Add10_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Add10_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No264_out_to_MUX_Add10_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add10_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Add10_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No114_out_to_Add23_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No115_out_to_Add23_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1043_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg725_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg915_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1046_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No183_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg607_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg483_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg483_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg984_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No116_out_to_Add23_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No117_out_to_Add23_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg919_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg945_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No118_out_to_Add23_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No119_out_to_Add23_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Add23_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out_to_MUX_Add23_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Add23_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Add23_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Add23_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out_to_MUX_Add23_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add23_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Add23_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Add23_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Add23_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Add23_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Add23_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out_to_MUX_Add23_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg990_out_to_MUX_Add23_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Add23_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out_to_MUX_Add23_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No185_out_to_MUX_Add23_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Add23_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add23_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add23_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out_to_MUX_Add23_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out_to_MUX_Add23_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out_to_MUX_Add23_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out_to_MUX_Add23_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No120_out_to_Add113_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No121_out_to_Add113_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out_to_MUX_Add113_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add113_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Add113_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add113_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Add113_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Add113_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Add113_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Add113_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Add113_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Add113_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1071_out_to_MUX_Add113_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No238_out_to_MUX_Add113_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out_to_MUX_Add113_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add113_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add113_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg604_out_to_MUX_Add113_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Add113_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out_to_MUX_Add113_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out_to_MUX_Add113_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Add113_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1004_out_to_MUX_Add113_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Add113_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1074_out_to_MUX_Add113_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg605_out_to_MUX_Add113_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No122_out_to_Add113_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No123_out_to_Add113_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Add113_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No239_out_to_MUX_Add113_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg483_out_to_MUX_Add113_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add113_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Add113_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out_to_MUX_Add113_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Add113_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Add113_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Add113_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out_to_MUX_Add113_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Add113_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg984_out_to_MUX_Add113_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out_to_MUX_Add113_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out_to_MUX_Add113_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Add113_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add113_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add113_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out_to_MUX_Add113_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg607_out_to_MUX_Add113_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out_to_MUX_Add113_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out_to_MUX_Add113_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg483_out_to_MUX_Add113_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out_to_MUX_Add113_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out_to_MUX_Add113_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No124_out_to_Add113_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No125_out_to_Add113_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out_to_MUX_Add113_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Add113_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1013_out_to_MUX_Add113_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Add113_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out_to_MUX_Add113_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add113_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Add113_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Add113_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Add113_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Add113_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Add113_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Add113_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Add113_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Add113_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1016_out_to_MUX_Add113_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No184_out_to_MUX_Add113_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Add113_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add113_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add113_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Add113_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Add113_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Add113_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Add113_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out_to_MUX_Add113_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No126_out_to_Add113_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No127_out_to_Add113_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Add113_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Add113_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Add113_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1018_out_to_MUX_Add113_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No241_out_to_MUX_Add113_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out_to_MUX_Add113_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add113_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Add113_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg731_out_to_MUX_Add113_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg731_out_to_MUX_Add113_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out_to_MUX_Add113_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out_to_MUX_Add113_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out_to_MUX_Add113_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Add113_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg756_out_to_MUX_Add113_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1021_out_to_MUX_Add113_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out_to_MUX_Add113_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Add113_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add113_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Add113_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out_to_MUX_Add113_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out_to_MUX_Add113_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Add113_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Add113_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No128_out_to_Add113_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No129_out_to_Add113_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Add113_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Add113_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out_to_MUX_Add113_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Add113_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Add113_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg994_out_to_MUX_Add113_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out_to_MUX_Add113_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Add113_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add113_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg408_out_to_MUX_Add113_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out_to_MUX_Add113_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out_to_MUX_Add113_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out_to_MUX_Add113_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out_to_MUX_Add113_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Add113_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Add113_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Add113_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_Add113_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No186_out_to_MUX_Add113_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out_to_MUX_Add113_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add113_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out_to_MUX_Add113_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg952_out_to_MUX_Add113_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Add113_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No130_out_to_Add24_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No131_out_to_Add24_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out_to_MUX_Add24_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Add24_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Add24_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Add24_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Add24_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out_to_MUX_Add24_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg736_out_to_MUX_Add24_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No221_out_to_MUX_Add24_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add24_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out_to_MUX_Add24_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg974_out_to_MUX_Add24_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out_to_MUX_Add24_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out_to_MUX_Add24_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg951_out_to_MUX_Add24_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out_to_MUX_Add24_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg951_out_to_MUX_Add24_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Add24_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Add24_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Add24_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No228_out_to_MUX_Add24_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add24_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Add24_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg930_out_to_MUX_Add24_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg952_out_to_MUX_Add24_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No132_out_to_Add32_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No133_out_to_Add32_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Add32_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Add32_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Add32_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Add32_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Add32_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Add32_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Add32_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1029_out_to_MUX_Add32_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out_to_MUX_Add32_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out_to_MUX_Add32_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Add32_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Add32_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg955_out_to_MUX_Add32_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out_to_MUX_Add32_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out_to_MUX_Add32_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out_to_MUX_Add32_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Add32_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Add32_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out_to_MUX_Add32_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1065_out_to_MUX_Add32_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No187_out_to_MUX_Add32_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out_to_MUX_Add32_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add32_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out_to_MUX_Add32_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No134_out_to_Add122_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No135_out_to_Add122_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No47_out_to_MUX_Add122_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Add122_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out_to_MUX_Add122_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Add122_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Add122_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out_to_MUX_Add122_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Add122_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Add122_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No243_out_to_MUX_Add122_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Add122_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add122_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out_to_MUX_Add122_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Add122_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Add122_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Add122_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out_to_MUX_Add122_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out_to_MUX_Add122_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out_to_MUX_Add122_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Add122_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Add122_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg620_out_to_MUX_Add122_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out_to_MUX_Add122_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add122_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Add122_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No136_out_to_Add33_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No137_out_to_Add33_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add33_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Add33_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Add33_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Add33_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add33_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add33_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add33_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Add33_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out_to_MUX_Add33_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1004_out_to_MUX_Add33_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Add33_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out_to_MUX_Add33_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out_to_MUX_Add33_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add33_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg721_out_to_MUX_Add33_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Add33_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg604_out_to_MUX_Add33_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out_to_MUX_Add33_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out_to_MUX_Add33_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out_to_MUX_Add33_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out_to_MUX_Add33_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Add33_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_Add33_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Add33_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No138_out_to_Add33_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No139_out_to_Add33_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg919_out_to_MUX_Add33_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Add33_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Add33_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No240_out_to_MUX_Add33_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out_to_MUX_Add33_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Add33_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Add33_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Add33_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Add33_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Add33_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Add33_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Add33_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg945_out_to_MUX_Add33_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg751_out_to_MUX_Add33_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Add33_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out_to_MUX_Add33_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out_to_MUX_Add33_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add33_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Add33_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg946_out_to_MUX_Add33_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Add33_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out_to_MUX_Add33_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out_to_MUX_Add33_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Add33_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No140_out_to_Add33_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No141_out_to_Add33_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Add33_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Add33_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Add33_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out_to_MUX_Add33_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Add33_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out_to_MUX_Add33_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No242_out_to_MUX_Add33_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Add33_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Add33_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out_to_MUX_Add33_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No46_out_to_MUX_Add33_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Add33_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg951_out_to_MUX_Add33_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out_to_MUX_Add33_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out_to_MUX_Add33_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out_to_MUX_Add33_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out_to_MUX_Add33_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Add33_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_Add33_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out_to_MUX_Add33_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add33_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Add33_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Add33_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out_to_MUX_Add33_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No142_out_to_Add33_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No143_out_to_Add33_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg977_out_to_MUX_Add33_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Add33_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Add33_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out_to_MUX_Add33_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Add33_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Add33_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_Add33_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out_to_MUX_Add33_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg740_out_to_MUX_Add33_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No222_out_to_MUX_Add33_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add33_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Add33_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Add33_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out_to_MUX_Add33_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg954_out_to_MUX_Add33_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Add33_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out_to_MUX_Add33_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg954_out_to_MUX_Add33_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Add33_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out_to_MUX_Add33_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Add33_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No229_out_to_MUX_Add33_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add33_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_Add33_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No144_out_to_Add33_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No145_out_to_Add33_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Add33_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out_to_MUX_Add33_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out_to_MUX_Add33_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Add33_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Add33_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out_to_MUX_Add33_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out_to_MUX_Add33_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1001_out_to_MUX_Add33_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1067_out_to_MUX_Add33_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out_to_MUX_Add33_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Add33_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Add33_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out_to_MUX_Add33_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out_to_MUX_Add33_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out_to_MUX_Add33_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out_to_MUX_Add33_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out_to_MUX_Add33_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out_to_MUX_Add33_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1033_out_to_MUX_Add33_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg601_out_to_MUX_Add33_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1080_out_to_MUX_Add33_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out_to_MUX_Add33_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out_to_MUX_Add33_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add33_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No146_out_to_Add123_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No147_out_to_Add123_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No217_out_to_MUX_Add123_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add123_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out_to_MUX_Add123_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Add123_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Add123_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out_to_MUX_Add123_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out_to_MUX_Add123_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add123_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Add123_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Add123_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out_to_MUX_Add123_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Add123_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No224_out_to_MUX_Add123_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add123_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Add123_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Add123_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Add123_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Add123_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Add123_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out_to_MUX_Add123_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Add123_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Add123_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out_to_MUX_Add123_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out_to_MUX_Add123_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No148_out_to_Add123_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No149_out_to_Add123_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out_to_MUX_Add123_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg724_out_to_MUX_Add123_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Add123_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Add123_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Add123_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Add123_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out_to_MUX_Add123_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Add123_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Add123_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Add123_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg915_out_to_MUX_Add123_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Add123_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Add123_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Add123_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out_to_MUX_Add123_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add123_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg725_out_to_MUX_Add123_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Add123_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out_to_MUX_Add123_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Add123_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Add123_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out_to_MUX_Add123_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Add123_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Add123_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No150_out_to_Add123_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No151_out_to_Add123_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Add123_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Add123_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Add123_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out_to_MUX_Add123_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Add123_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add123_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg536_out_to_MUX_Add123_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No44_out_to_MUX_Add123_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out_to_MUX_Add123_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg919_out_to_MUX_Add123_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg919_out_to_MUX_Add123_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Add123_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg946_out_to_MUX_Add123_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Add123_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Add123_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out_to_MUX_Add123_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Add123_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add123_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out_to_MUX_Add123_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out_to_MUX_Add123_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Add123_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg945_out_to_MUX_Add123_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg945_out_to_MUX_Add123_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out_to_MUX_Add123_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No152_out_to_Add123_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No153_out_to_Add123_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out_to_MUX_Add123_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg923_out_to_MUX_Add123_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Add123_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Add123_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out_to_MUX_Add123_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Add123_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Add123_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Add123_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out_to_MUX_Add123_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out_to_MUX_Add123_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg923_out_to_MUX_Add123_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg923_out_to_MUX_Add123_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Add123_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Add123_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Add123_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Add123_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out_to_MUX_Add123_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out_to_MUX_Add123_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add123_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out_to_MUX_Add123_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg949_out_to_MUX_Add123_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Add123_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Add123_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Add123_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No154_out_to_Add123_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No155_out_to_Add123_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out_to_MUX_Add123_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out_to_MUX_Add123_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out_to_MUX_Add123_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_Add123_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_Add123_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Add123_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Add123_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Add123_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out_to_MUX_Add123_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Add123_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No223_out_to_MUX_Add123_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add123_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out_to_MUX_Add123_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg958_out_to_MUX_Add123_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out_to_MUX_Add123_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Add123_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Add123_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out_to_MUX_Add123_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add123_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out_to_MUX_Add123_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Add123_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Add123_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No230_out_to_MUX_Add123_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add123_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No156_out_to_Add35_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No157_out_to_Add35_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Add35_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add35_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg823_out_to_MUX_Add35_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No42_out_to_MUX_Add35_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out_to_MUX_Add35_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Add35_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Add35_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out_to_MUX_Add35_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Add35_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_Add35_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg626_out_to_MUX_Add35_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg961_out_to_MUX_Add35_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No259_out_to_MUX_Add35_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add35_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out_to_MUX_Add35_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Add35_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg481_out_to_MUX_Add35_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Add35_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Add35_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Add35_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Add35_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1041_out_to_MUX_Add35_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Add35_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Add35_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No158_out_to_Add35_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No159_out_to_Add35_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg629_out_to_MUX_Add35_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg915_out_to_MUX_Add35_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No218_out_to_MUX_Add35_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add35_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg533_out_to_MUX_Add35_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No43_out_to_MUX_Add35_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Add35_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg915_out_to_MUX_Add35_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg915_out_to_MUX_Add35_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Add35_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Add35_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1007_out_to_MUX_Add35_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Add35_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out_to_MUX_Add35_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No225_out_to_MUX_Add35_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add35_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Add35_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Add35_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Add35_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Add35_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Add35_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Add35_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Add35_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out_to_MUX_Add35_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No160_out_to_Add35_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No161_out_to_Add35_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out_to_MUX_Add35_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No48_out_to_MUX_Add35_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out_to_MUX_Add35_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Add35_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Add35_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_Add35_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Add35_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1033_out_to_MUX_Add35_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Add35_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg979_out_to_MUX_Add35_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Add35_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add35_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out_to_MUX_Add35_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Add35_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg958_out_to_MUX_Add35_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_Add35_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_Add35_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Add35_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_Add35_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1069_out_to_MUX_Add35_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_Add35_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_Add35_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No265_out_to_MUX_Add35_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add35_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No162_out_to_Add130_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No163_out_to_Add130_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add130_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg644_out_to_MUX_Add130_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out_to_MUX_Add130_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg980_out_to_MUX_Add130_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add130_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Add130_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg958_out_to_MUX_Add130_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Add130_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No164_out_to_Product4_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No165_out_to_Product4_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg982_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1143_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1133_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1072_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No166_out_to_Product4_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No167_out_to_Product4_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg985_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1143_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1133_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1083_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No168_out_to_Product4_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No169_out_to_Product4_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1143_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1133_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1049_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No170_out_to_Product4_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No171_out_to_Product4_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1143_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1133_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1055_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No172_out_to_Product4_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No173_out_to_Product4_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg690_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1143_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1133_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1023_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No174_out_to_Product4_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No175_out_to_Product4_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1143_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1133_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1030_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No176_out_to_Product4_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No177_out_to_Product4_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1143_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1133_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1068_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No178_out_to_Product21_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No179_out_to_Product21_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1132_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1072_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1039_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1145_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No180_out_to_Product21_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No181_out_to_Product21_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1132_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1083_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1044_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1145_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No182_out_to_Product21_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No183_out_to_Product21_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1132_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1049_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1014_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1145_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No184_out_to_Product21_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No185_out_to_Product21_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1132_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1055_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1055_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1145_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No186_out_to_Product21_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No187_out_to_Product21_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1132_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1023_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1023_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1145_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No188_out_to_Product21_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No189_out_to_Product21_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1132_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1030_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg999_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1145_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No190_out_to_Product21_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No191_out_to_Product21_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1132_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1068_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1068_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1145_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No192_out_to_Subtract2_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No193_out_to_Subtract2_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg604_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No7_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No194_out_to_Subtract2_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No195_out_to_Subtract2_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg963_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No196_out_to_Subtract2_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No197_out_to_Subtract2_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg892_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg536_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1014_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg967_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No198_out_to_Subtract2_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No199_out_to_Subtract2_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg895_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1019_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg969_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg757_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No200_out_to_Subtract2_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No201_out_to_Subtract2_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1023_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg408_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg972_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg972_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg706_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg972_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No202_out_to_Subtract2_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No203_out_to_Subtract2_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg765_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg975_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No204_out_to_Subtract2_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No205_out_to_Subtract2_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg500_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No13_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No206_out_to_Product5_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No207_out_to_Product5_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1127_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1132_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1147_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1004_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg982_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1096_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No208_out_to_Product5_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No209_out_to_Product5_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1127_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1132_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1147_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1007_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg985_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No210_out_to_Product5_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No211_out_to_Product5_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1132_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1147_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1127_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg878_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg986_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No212_out_to_Product5_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No213_out_to_Product5_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1132_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1147_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1127_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1017_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No214_out_to_Product5_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No215_out_to_Product5_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1127_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1132_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1147_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg993_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg690_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No216_out_to_Product5_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No217_out_to_Product5_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out_to_MUX_Product5_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product5_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product5_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1127_out_to_MUX_Product5_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Product5_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1132_out_to_MUX_Product5_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1147_out_to_MUX_Product5_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product5_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product5_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product5_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product5_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out_to_MUX_Product5_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Product5_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Product5_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product5_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_Product5_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Product5_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Product5_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1061_out_to_MUX_Product5_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_Product5_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product5_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Product5_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Product5_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Product5_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No218_out_to_Product5_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No219_out_to_Product5_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out_to_MUX_Product5_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out_to_MUX_Product5_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product5_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product5_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1127_out_to_MUX_Product5_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Product5_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1132_out_to_MUX_Product5_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1147_out_to_MUX_Product5_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product5_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product5_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product5_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product5_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Product5_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Product5_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Product5_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Product5_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1033_out_to_MUX_Product5_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product5_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out_to_MUX_Product5_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1077_out_to_MUX_Product5_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product5_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product5_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product5_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Product5_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No220_out_to_Product12_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No221_out_to_Product12_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1146_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1133_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1151_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1094_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1039_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1096_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No222_out_to_Product12_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No223_out_to_Product12_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1146_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1133_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1151_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1044_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No224_out_to_Product12_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No225_out_to_Product12_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1133_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1151_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1146_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1014_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg878_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No226_out_to_Product12_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No227_out_to_Product12_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1133_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1151_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1146_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1055_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No228_out_to_Product12_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No229_out_to_Product12_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1146_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1133_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1151_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1023_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No230_out_to_Product12_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No231_out_to_Product12_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Product12_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product12_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Product12_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1146_out_to_MUX_Product12_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Product12_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1133_out_to_MUX_Product12_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1151_out_to_MUX_Product12_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Product12_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product12_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Product12_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Product12_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Product12_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out_to_MUX_Product12_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product12_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product12_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1060_out_to_MUX_Product12_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Product12_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg999_out_to_MUX_Product12_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1061_out_to_MUX_Product12_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product12_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product12_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product12_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product12_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out_to_MUX_Product12_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No232_out_to_Product12_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No233_out_to_Product12_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Product12_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Product12_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product12_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product12_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1146_out_to_MUX_Product12_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Product12_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1133_out_to_MUX_Product12_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1151_out_to_MUX_Product12_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Product12_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product12_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Product12_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product12_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out_to_MUX_Product12_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out_to_MUX_Product12_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product12_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product12_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1088_out_to_MUX_Product12_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product12_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1068_out_to_MUX_Product12_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1077_out_to_MUX_Product12_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product12_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product12_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product12_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product12_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No234_out_to_Product22_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No235_out_to_Product22_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1094_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1150_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1005_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No236_out_to_Product22_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No237_out_to_Product22_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1150_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1008_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No238_out_to_Product22_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No239_out_to_Product22_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg987_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1150_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No240_out_to_Product22_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No241_out_to_Product22_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg991_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1150_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No242_out_to_Product22_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No243_out_to_Product22_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1150_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No244_out_to_Product22_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No245_out_to_Product22_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product22_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out_to_MUX_Product22_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product22_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1060_out_to_MUX_Product22_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Product22_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_Product22_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product22_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product22_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product22_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Product22_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product22_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product22_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Product22_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Product22_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Product22_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1150_out_to_MUX_Product22_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Product22_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg869_out_to_MUX_Product22_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product22_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Product22_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Product22_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Product22_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Product22_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Product22_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No246_out_to_Product22_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No247_out_to_Product22_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product22_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product22_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out_to_MUX_Product22_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product22_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1088_out_to_MUX_Product22_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Product22_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_Product22_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product22_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product22_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product22_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Product22_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product22_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Product22_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Product22_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Product22_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Product22_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1150_out_to_MUX_Product22_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product22_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1002_out_to_MUX_Product22_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product22_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Product22_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Product22_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Product22_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Product22_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No248_out_to_Product32_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No249_out_to_Product32_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1154_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg666_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg775_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1038_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No250_out_to_Product32_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No251_out_to_Product32_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1154_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1043_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No252_out_to_Product32_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No253_out_to_Product32_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1154_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1013_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No254_out_to_Product32_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No255_out_to_Product32_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1154_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1018_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg705_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No256_out_to_Product32_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No257_out_to_Product32_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1154_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg994_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No258_out_to_Product32_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No259_out_to_Product32_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1154_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No260_out_to_Product32_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No261_out_to_Product32_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1154_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1101_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1034_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No262_out_to_Subtract3_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No263_out_to_Subtract3_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg960_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg667_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No264_out_to_Subtract3_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No265_out_to_Subtract3_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg483_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg724_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg533_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1009_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg964_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No266_out_to_Subtract3_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No267_out_to_Subtract3_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg891_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg891_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg986_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg966_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg966_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No268_out_to_Subtract3_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No269_out_to_Subtract3_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg896_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg877_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg895_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg895_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg970_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg634_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg969_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg969_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No270_out_to_Subtract3_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No271_out_to_Subtract3_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg993_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg705_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No214_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg952_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg973_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg953_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg973_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No272_out_to_Subtract3_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No273_out_to_Subtract3_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Subtract3_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Subtract3_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Subtract3_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1030_out_to_MUX_Subtract3_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out_to_MUX_Subtract3_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Subtract3_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out_to_MUX_Subtract3_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Subtract3_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out_to_MUX_Subtract3_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No215_out_to_MUX_Subtract3_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract3_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg955_out_to_MUX_Subtract3_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg976_out_to_MUX_Subtract3_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg975_out_to_MUX_Subtract3_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg975_out_to_MUX_Subtract3_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Subtract3_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Subtract3_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg976_out_to_MUX_Subtract3_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Subtract3_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Subtract3_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Subtract3_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out_to_MUX_Subtract3_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract3_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg956_out_to_MUX_Subtract3_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No274_out_to_Subtract3_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No275_out_to_Subtract3_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No276_out_to_Product6_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No277_out_to_Product6_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg775_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1128_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1138_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1156_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg982_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1005_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No278_out_to_Product6_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No279_out_to_Product6_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1128_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1138_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1156_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg985_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1008_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No280_out_to_Product6_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No281_out_to_Product6_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1138_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1128_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg987_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1156_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No282_out_to_Product6_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No283_out_to_Product6_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1128_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1138_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg705_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg991_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg991_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1156_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No284_out_to_Product6_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No285_out_to_Product6_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1128_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1138_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1156_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No286_out_to_Product6_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No287_out_to_Product6_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out_to_MUX_Product6_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product6_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product6_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_Product6_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1128_out_to_MUX_Product6_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1138_out_to_MUX_Product6_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product6_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product6_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product6_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product6_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product6_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Product6_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Product6_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Product6_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Product6_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1156_out_to_MUX_Product6_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Product6_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg869_out_to_MUX_Product6_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Product6_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Product6_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Product6_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Product6_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Product6_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Product6_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No288_out_to_Product6_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No289_out_to_Product6_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Product6_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out_to_MUX_Product6_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product6_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product6_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1101_out_to_MUX_Product6_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1128_out_to_MUX_Product6_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1138_out_to_MUX_Product6_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product6_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product6_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product6_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product6_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product6_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Product6_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Product6_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product6_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Product6_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1156_out_to_MUX_Product6_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1002_out_to_MUX_Product6_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1002_out_to_MUX_Product6_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Product6_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Product6_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Product6_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Product6_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Product6_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No290_out_to_Product23_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No291_out_to_Product23_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg666_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1130_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1038_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg982_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1138_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No292_out_to_Product23_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No293_out_to_Product23_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1130_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1043_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg985_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1138_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No294_out_to_Product23_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No295_out_to_Product23_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1013_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1130_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1138_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No296_out_to_Product23_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No297_out_to_Product23_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1130_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1018_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg991_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1138_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No298_out_to_Product23_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No299_out_to_Product23_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1130_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg994_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1138_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No300_out_to_Product23_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No301_out_to_Product23_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Product23_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product23_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Product23_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Product23_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1130_out_to_MUX_Product23_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_Product23_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product23_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Product23_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Product23_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Product23_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Product23_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Product23_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out_to_MUX_Product23_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Product23_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product23_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Product23_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Product23_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1138_out_to_MUX_Product23_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Product23_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product23_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product23_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product23_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product23_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Product23_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No302_out_to_Product23_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No303_out_to_Product23_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Product23_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product23_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product23_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product23_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Product23_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1130_out_to_MUX_Product23_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1034_out_to_MUX_Product23_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product23_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Product23_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product23_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Product23_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product23_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Product23_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out_to_MUX_Product23_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Product23_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product23_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product23_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1002_out_to_MUX_Product23_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1138_out_to_MUX_Product23_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Product23_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product23_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product23_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product23_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product23_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No304_out_to_Product33_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No305_out_to_Product33_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1005_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1142_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg981_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1094_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1099_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1130_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1072_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg981_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1073_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No306_out_to_Product33_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No307_out_to_Product33_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1008_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1142_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1045_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1081_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1130_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1083_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No308_out_to_Product33_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No309_out_to_Product33_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1142_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg987_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1049_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1015_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1047_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1052_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1130_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No310_out_to_Product33_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No311_out_to_Product33_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1018_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1142_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1130_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1056_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1058_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No312_out_to_Product33_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No313_out_to_Product33_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg994_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1142_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1025_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1130_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg995_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No314_out_to_Product33_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No315_out_to_Product33_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg869_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1142_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1130_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1030_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1000_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No316_out_to_Product33_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No317_out_to_Product33_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1034_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1142_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1001_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1003_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1093_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1130_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1077_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1001_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1078_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1001_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1101_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No318_out_to_Subtract4_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No319_out_to_Subtract4_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No210_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg646_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1006_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg961_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No320_out_to_Subtract4_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No321_out_to_Subtract4_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No211_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg649_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg649_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg508_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg963_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg963_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1007_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No322_out_to_Subtract4_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No323_out_to_Subtract4_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No212_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg946_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg892_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg536_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1012_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1049_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg879_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg512_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg967_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No324_out_to_Subtract4_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No325_out_to_Subtract4_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No213_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg949_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1017_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1055_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1017_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg950_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg634_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No326_out_to_Subtract4_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No327_out_to_Subtract4_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg705_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg463_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No270_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No328_out_to_Subtract4_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No329_out_to_Subtract4_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg620_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg997_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No271_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No330_out_to_Subtract4_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No331_out_to_Subtract4_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg958_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1035_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg771_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No216_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg959_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg978_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg602_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg978_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg528_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No332_out_to_Subtract5_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No333_out_to_Subtract5_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg616_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg736_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No334_out_to_Subtract5_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No335_out_to_Subtract5_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out_to_MUX_Subtract5_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out_to_MUX_Subtract5_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out_to_MUX_Subtract5_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract5_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract5_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out_to_MUX_Subtract5_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Subtract5_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out_to_MUX_Subtract5_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Subtract5_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Subtract5_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract5_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg740_out_to_MUX_Subtract5_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_Subtract5_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out_to_MUX_Subtract5_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out_to_MUX_Subtract5_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out_to_MUX_Subtract5_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out_to_MUX_Subtract5_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Subtract5_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Subtract5_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Subtract5_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract5_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract5_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract5_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Subtract5_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No336_out_to_Product26_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No337_out_to_Product26_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1144_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1105_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1004_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1038_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg981_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg983_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1098_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1071_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1004_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1097_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No338_out_to_Product26_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No339_out_to_Product26_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1144_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1105_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg984_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1084_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg984_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1008_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1085_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1082_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No340_out_to_Product26_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No341_out_to_Product26_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1105_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1144_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1050_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg987_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg680_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1051_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1048_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No342_out_to_Product26_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No343_out_to_Product26_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1144_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1105_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg991_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg990_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No344_out_to_Product26_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No345_out_to_Product26_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1144_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1105_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1024_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg994_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No346_out_to_Product26_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No347_out_to_Product26_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product26_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product26_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product26_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product26_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1144_out_to_MUX_Product26_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1105_out_to_MUX_Product26_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product26_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product26_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product26_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product26_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product26_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product26_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_Product26_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg870_out_to_MUX_Product26_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg774_out_to_MUX_Product26_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Product26_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1029_out_to_MUX_Product26_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Product26_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Product26_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_Product26_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1031_out_to_MUX_Product26_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg997_out_to_MUX_Product26_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1029_out_to_MUX_Product26_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Product26_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No348_out_to_Product26_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No349_out_to_Product26_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product26_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product26_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product26_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product26_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product26_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1144_out_to_MUX_Product26_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1105_out_to_MUX_Product26_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product26_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product26_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product26_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product26_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product26_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Product26_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1033_out_to_MUX_Product26_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1036_out_to_MUX_Product26_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1092_out_to_MUX_Product26_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product26_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out_to_MUX_Product26_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Product26_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Product26_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1033_out_to_MUX_Product26_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1091_out_to_MUX_Product26_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1033_out_to_MUX_Product26_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1067_out_to_MUX_Product26_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No350_out_to_Subtract7_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No351_out_to_Subtract7_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg891_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg966_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg510_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No352_out_to_Subtract7_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No353_out_to_Subtract7_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No10_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No354_out_to_Subtract7_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No355_out_to_Subtract7_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg864_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg408_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No356_out_to_Subtract7_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No357_out_to_Subtract7_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Subtract7_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract7_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract7_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Subtract7_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Subtract7_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out_to_MUX_Subtract7_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg952_out_to_MUX_Subtract7_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Subtract7_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract7_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract7_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract7_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out_to_MUX_Subtract7_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out_to_MUX_Subtract7_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out_to_MUX_Subtract7_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out_to_MUX_Subtract7_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Subtract7_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Subtract7_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Subtract7_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg972_out_to_MUX_Subtract7_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg588_out_to_MUX_Subtract7_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract7_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract7_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract7_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Subtract7_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No358_out_to_Subtract7_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No359_out_to_Subtract7_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out_to_MUX_Subtract7_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg470_out_to_MUX_Subtract7_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out_to_MUX_Subtract7_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Subtract7_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Subtract7_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Subtract7_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_Subtract7_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Subtract7_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg955_out_to_MUX_Subtract7_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out_to_MUX_Subtract7_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Subtract7_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract7_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out_to_MUX_Subtract7_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out_to_MUX_Subtract7_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Subtract7_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Subtract7_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Subtract7_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Subtract7_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Subtract7_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Subtract7_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg975_out_to_MUX_Subtract7_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Subtract7_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract7_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract7_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No360_out_to_Subtract8_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No361_out_to_Subtract8_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Subtract8_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Subtract8_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract8_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Subtract8_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Subtract8_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg485_out_to_MUX_Subtract8_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Subtract8_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Subtract8_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Subtract8_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Subtract8_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg483_out_to_MUX_Subtract8_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg607_out_to_MUX_Subtract8_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Subtract8_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract8_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract8_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out_to_MUX_Subtract8_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Subtract8_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No8_out_to_MUX_Subtract8_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Subtract8_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Subtract8_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Subtract8_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Subtract8_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Subtract8_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Subtract8_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No362_out_to_Subtract8_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No363_out_to_Subtract8_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No9_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No364_out_to_Subtract8_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No365_out_to_Subtract8_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1018_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg949_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg688_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg990_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1021_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg969_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No11_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No366_out_to_Subtract8_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No367_out_to_Subtract8_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out_to_MUX_Subtract8_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Subtract8_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Subtract8_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Subtract8_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Subtract8_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg994_out_to_MUX_Subtract8_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out_to_MUX_Subtract8_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Subtract8_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract8_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract8_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Subtract8_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out_to_MUX_Subtract8_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No12_out_to_MUX_Subtract8_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Subtract8_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_Subtract8_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Subtract8_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out_to_MUX_Subtract8_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_Subtract8_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out_to_MUX_Subtract8_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Subtract8_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract8_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract8_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Subtract8_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out_to_MUX_Subtract8_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No368_out_to_Product18_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No369_out_to_Product18_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1155_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg981_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1094_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1099_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg775_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg981_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1073_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No370_out_to_Product18_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No371_out_to_Product18_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1155_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1045_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1081_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No372_out_to_Product18_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No373_out_to_Product18_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1155_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1015_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1047_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1052_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No374_out_to_Product18_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No375_out_to_Product18_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1155_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1056_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1058_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No376_out_to_Product18_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No377_out_to_Product18_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1155_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1025_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg995_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No378_out_to_Product18_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No379_out_to_Product18_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Product18_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Product18_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product18_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Product18_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1155_out_to_MUX_Product18_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Product18_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product18_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product18_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product18_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Product18_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product18_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out_to_MUX_Product18_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Product18_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out_to_MUX_Product18_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out_to_MUX_Product18_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product18_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_Product18_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Product18_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Product18_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Product18_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1000_out_to_MUX_Product18_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_Product18_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_Product18_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Product18_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No380_out_to_Product18_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No381_out_to_Product18_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out_to_MUX_Product18_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Product18_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Product18_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product18_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Product18_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1155_out_to_MUX_Product18_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Product18_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product18_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product18_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product18_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Product18_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product18_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product18_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1001_out_to_MUX_Product18_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1003_out_to_MUX_Product18_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1093_out_to_MUX_Product18_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product18_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1088_out_to_MUX_Product18_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Product18_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Product18_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1001_out_to_MUX_Product18_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1078_out_to_MUX_Product18_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1001_out_to_MUX_Product18_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1101_out_to_MUX_Product18_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No382_out_to_Product28_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No383_out_to_Product28_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1004_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1038_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg981_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg983_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1098_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1157_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1105_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1004_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1097_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg775_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No384_out_to_Product28_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No385_out_to_Product28_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg984_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1084_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg984_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1008_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1085_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1157_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1105_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No386_out_to_Product28_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No387_out_to_Product28_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1105_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1050_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg987_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg680_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1051_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1157_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No388_out_to_Product28_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No389_out_to_Product28_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1157_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1105_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg991_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg990_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No390_out_to_Product28_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No391_out_to_Product28_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1157_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1105_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1024_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg994_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No392_out_to_Product28_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No393_out_to_Product28_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_Product28_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg870_out_to_MUX_Product28_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg774_out_to_MUX_Product28_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Product28_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1157_out_to_MUX_Product28_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1105_out_to_MUX_Product28_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Product28_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_Product28_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1031_out_to_MUX_Product28_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg997_out_to_MUX_Product28_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1029_out_to_MUX_Product28_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Product28_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Product28_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Product28_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product28_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Product28_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_Product28_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Product28_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product28_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product28_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product28_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Product28_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product28_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out_to_MUX_Product28_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No394_out_to_Product28_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No395_out_to_Product28_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1033_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1036_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1092_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1157_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1105_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1033_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1091_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1033_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1067_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1088_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No396_out_to_Subtract9_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No397_out_to_Subtract9_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg646_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg434_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg666_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No266_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg960_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg960_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg982_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg604_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No398_out_to_Subtract9_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No399_out_to_Subtract9_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg890_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg533_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1007_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1044_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1084_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg607_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No267_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg944_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg964_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No400_out_to_Subtract9_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No401_out_to_Subtract9_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg894_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No268_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg894_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No402_out_to_Subtract9_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No403_out_to_Subtract9_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg898_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg896_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No269_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg970_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No404_out_to_Subtract9_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No405_out_to_Subtract9_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg705_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg408_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg616_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No46_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No406_out_to_Subtract9_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No407_out_to_Subtract9_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg905_out_to_MUX_Subtract9_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_Subtract9_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Subtract9_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1061_out_to_MUX_Subtract9_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Subtract9_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Subtract9_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out_to_MUX_Subtract9_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Subtract9_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Subtract9_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out_to_MUX_Subtract9_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Subtract9_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract9_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No47_out_to_MUX_Subtract9_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Subtract9_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Subtract9_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_Subtract9_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out_to_MUX_Subtract9_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Subtract9_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out_to_MUX_Subtract9_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Subtract9_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out_to_MUX_Subtract9_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Subtract9_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract9_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract9_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No408_out_to_Subtract9_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No409_out_to_Subtract9_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract9_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out_to_MUX_Subtract9_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Subtract9_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Subtract9_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Subtract9_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Subtract9_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Subtract9_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Subtract9_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Subtract9_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Subtract9_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Subtract9_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract9_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Subtract9_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out_to_MUX_Subtract9_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out_to_MUX_Subtract9_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg978_out_to_MUX_Subtract9_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Subtract9_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Subtract9_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg979_out_to_MUX_Subtract9_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1002_out_to_MUX_Subtract9_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Subtract9_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out_to_MUX_Subtract9_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No272_out_to_MUX_Subtract9_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract9_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No410_out_to_Subtract10_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No411_out_to_Subtract10_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg946_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg966_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No412_out_to_Product50_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No413_out_to_Product50_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1149_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1148_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1070_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1040_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1100_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No414_out_to_Product50_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No415_out_to_Product50_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1148_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1149_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1007_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1042_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1010_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1087_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No416_out_to_Product50_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No417_out_to_Product50_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1148_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1149_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg986_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg878_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1012_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg988_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1053_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No418_out_to_Product50_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No419_out_to_Product50_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1148_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1149_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg990_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1017_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1020_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1059_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No420_out_to_Product50_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No421_out_to_Product50_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1148_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1149_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1026_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg705_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1022_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1024_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No422_out_to_Product50_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No423_out_to_Product50_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product50_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product50_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product50_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product50_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Product50_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Product50_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product50_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1148_out_to_MUX_Product50_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product50_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product50_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1149_out_to_MUX_Product50_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product50_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out_to_MUX_Product50_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1031_out_to_MUX_Product50_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1064_out_to_MUX_Product50_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out_to_MUX_Product50_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Product50_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Product50_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product50_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg997_out_to_MUX_Product50_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out_to_MUX_Product50_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1060_out_to_MUX_Product50_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Product50_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_Product50_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No424_out_to_Product50_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No425_out_to_Product50_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product50_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product50_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product50_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product50_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product50_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out_to_MUX_Product50_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product50_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product50_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1148_out_to_MUX_Product50_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product50_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product50_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1149_out_to_MUX_Product50_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out_to_MUX_Product50_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Product50_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1078_out_to_MUX_Product50_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1079_out_to_MUX_Product50_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Product50_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Product50_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Product50_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out_to_MUX_Product50_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1066_out_to_MUX_Product50_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1090_out_to_MUX_Product50_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1075_out_to_MUX_Product50_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out_to_MUX_Product50_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No426_out_to_Product122_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No427_out_to_Product122_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1149_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1148_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1094_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1004_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg981_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg666_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1073_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1095_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1070_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No428_out_to_Product122_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No429_out_to_Product122_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1148_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1149_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1042_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1081_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg984_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1045_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No430_out_to_Product122_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No431_out_to_Product122_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1148_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1149_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1012_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg879_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1047_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1015_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No432_out_to_Product122_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No433_out_to_Product122_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1148_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1149_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1017_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1054_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg990_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1056_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No434_out_to_Product122_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No435_out_to_Product122_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1148_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1149_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg993_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg993_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No436_out_to_Product122_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No437_out_to_Product122_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product122_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product122_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product122_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out_to_MUX_Product122_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Product122_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Product122_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product122_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1148_out_to_MUX_Product122_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product122_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product122_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1149_out_to_MUX_Product122_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product122_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Product122_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1062_out_to_MUX_Product122_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out_to_MUX_Product122_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product122_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Product122_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Product122_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product122_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1028_out_to_MUX_Product122_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1062_out_to_MUX_Product122_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_Product122_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg997_out_to_MUX_Product122_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg997_out_to_MUX_Product122_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No438_out_to_Product122_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No439_out_to_Product122_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product122_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product122_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product122_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product122_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Product122_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Product122_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Product122_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product122_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1148_out_to_MUX_Product122_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product122_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product122_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1149_out_to_MUX_Product122_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1001_out_to_MUX_Product122_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out_to_MUX_Product122_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1091_out_to_MUX_Product122_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1089_out_to_MUX_Product122_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product122_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out_to_MUX_Product122_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Product122_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out_to_MUX_Product122_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1075_out_to_MUX_Product122_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1102_out_to_MUX_Product122_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1088_out_to_MUX_Product122_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1066_out_to_MUX_Product122_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No440_out_to_Product221_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No441_out_to_Product221_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1153_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1159_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1070_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1040_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1100_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg666_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg667_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No442_out_to_Product221_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No443_out_to_Product221_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1153_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1159_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1007_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1042_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1010_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1087_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No444_out_to_Product221_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No445_out_to_Product221_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1153_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1159_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg986_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg878_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1012_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg988_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1053_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No446_out_to_Product221_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No447_out_to_Product221_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1159_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1153_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg990_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1017_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1020_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1059_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No448_out_to_Product221_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No449_out_to_Product221_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1159_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1153_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1026_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1022_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1024_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No450_out_to_Product221_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No451_out_to_Product221_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Product221_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Product221_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product221_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_Product221_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1159_out_to_MUX_Product221_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out_to_MUX_Product221_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product221_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out_to_MUX_Product221_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product221_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Product221_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1153_out_to_MUX_Product221_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Product221_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out_to_MUX_Product221_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1031_out_to_MUX_Product221_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1064_out_to_MUX_Product221_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out_to_MUX_Product221_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg465_out_to_MUX_Product221_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Product221_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Product221_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg997_out_to_MUX_Product221_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out_to_MUX_Product221_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1060_out_to_MUX_Product221_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Product221_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_Product221_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No452_out_to_Product221_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No453_out_to_Product221_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Product221_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Product221_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Product221_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product221_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_Product221_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1159_out_to_MUX_Product221_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product221_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product221_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out_to_MUX_Product221_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product221_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Product221_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1153_out_to_MUX_Product221_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out_to_MUX_Product221_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Product221_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1078_out_to_MUX_Product221_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1079_out_to_MUX_Product221_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Product221_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Product221_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Product221_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Product221_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1066_out_to_MUX_Product221_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1090_out_to_MUX_Product221_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1075_out_to_MUX_Product221_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out_to_MUX_Product221_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No454_out_to_Product321_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No455_out_to_Product321_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1094_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1004_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg981_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg666_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1073_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1095_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1105_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1070_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1153_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1159_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No456_out_to_Product321_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No457_out_to_Product321_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1042_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1081_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg984_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1045_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1105_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1153_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1159_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No458_out_to_Product321_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No459_out_to_Product321_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1105_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1012_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg879_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1047_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1015_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1153_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1159_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No460_out_to_Product321_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No461_out_to_Product321_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1105_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1017_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1054_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg990_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1056_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1159_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1153_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No462_out_to_Product321_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No463_out_to_Product321_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg690_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1105_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg993_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg993_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1159_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1153_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No464_out_to_Product321_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No465_out_to_Product321_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Product321_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1062_out_to_MUX_Product321_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out_to_MUX_Product321_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_Product321_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out_to_MUX_Product321_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1105_out_to_MUX_Product321_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product321_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1028_out_to_MUX_Product321_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1062_out_to_MUX_Product321_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_Product321_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg997_out_to_MUX_Product321_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg997_out_to_MUX_Product321_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Product321_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Product321_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product321_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Product321_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1159_out_to_MUX_Product321_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Product321_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Product321_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out_to_MUX_Product321_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product321_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Product321_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1153_out_to_MUX_Product321_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Product321_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No466_out_to_Product321_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No467_out_to_Product321_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1001_out_to_MUX_Product321_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out_to_MUX_Product321_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1091_out_to_MUX_Product321_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1089_out_to_MUX_Product321_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_Product321_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out_to_MUX_Product321_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1105_out_to_MUX_Product321_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Product321_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1075_out_to_MUX_Product321_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1102_out_to_MUX_Product321_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1088_out_to_MUX_Product321_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1066_out_to_MUX_Product321_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Product321_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Product321_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Product321_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Product321_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out_to_MUX_Product321_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1159_out_to_MUX_Product321_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out_to_MUX_Product321_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product321_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out_to_MUX_Product321_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product321_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Product321_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1153_out_to_MUX_Product321_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No468_out_to_Subtract23_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No469_out_to_Subtract23_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1004_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1039_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1073_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No168_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg961_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg670_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No470_out_to_Subtract23_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No471_out_to_Subtract23_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1008_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No169_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg649_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No15_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg890_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No472_out_to_Subtract23_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No473_out_to_Subtract23_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg681_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg987_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No170_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg893_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No16_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No44_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg510_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No474_out_to_Subtract23_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No475_out_to_Subtract23_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Subtract23_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Subtract23_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Subtract23_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Subtract23_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No171_out_to_MUX_Subtract23_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out_to_MUX_Subtract23_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract23_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract23_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out_to_MUX_Subtract23_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Subtract23_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Subtract23_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Subtract23_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Subtract23_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Subtract23_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg881_out_to_MUX_Subtract23_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Subtract23_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Subtract23_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Subtract23_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract23_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract23_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg898_out_to_MUX_Subtract23_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Subtract23_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Subtract23_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Subtract23_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No476_out_to_Subtract23_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No477_out_to_Subtract23_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Subtract23_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out_to_MUX_Subtract23_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Subtract23_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Subtract23_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out_to_MUX_Subtract23_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out_to_MUX_Subtract23_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No172_out_to_MUX_Subtract23_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg972_out_to_MUX_Subtract23_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Subtract23_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract23_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg761_out_to_MUX_Subtract23_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Subtract23_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out_to_MUX_Subtract23_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Subtract23_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out_to_MUX_Subtract23_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out_to_MUX_Subtract23_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg762_out_to_MUX_Subtract23_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No18_out_to_MUX_Subtract23_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_Subtract23_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Subtract23_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract23_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract23_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Subtract23_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg973_out_to_MUX_Subtract23_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No478_out_to_Subtract23_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No479_out_to_Subtract23_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out_to_MUX_Subtract23_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Subtract23_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out_to_MUX_Subtract23_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Subtract23_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Subtract23_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Subtract23_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Subtract23_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_Subtract23_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No173_out_to_MUX_Subtract23_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg975_out_to_MUX_Subtract23_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract23_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract23_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out_to_MUX_Subtract23_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out_to_MUX_Subtract23_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg869_out_to_MUX_Subtract23_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Subtract23_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Subtract23_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Subtract23_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Subtract23_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No19_out_to_MUX_Subtract23_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg844_out_to_MUX_Subtract23_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Subtract23_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract23_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract23_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No480_out_to_Subtract23_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No481_out_to_Subtract23_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract23_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Subtract23_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out_to_MUX_Subtract23_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1033_out_to_MUX_Subtract23_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1068_out_to_MUX_Subtract23_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1078_out_to_MUX_Subtract23_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out_to_MUX_Subtract23_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Subtract23_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Subtract23_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No174_out_to_MUX_Subtract23_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Subtract23_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract23_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract23_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg979_out_to_MUX_Subtract23_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out_to_MUX_Subtract23_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Subtract23_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out_to_MUX_Subtract23_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_Subtract23_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1066_out_to_MUX_Subtract23_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Subtract23_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out_to_MUX_Subtract23_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out_to_MUX_Subtract23_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out_to_MUX_Subtract23_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract23_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No482_out_to_Subtract30_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No483_out_to_Subtract30_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg960_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg605_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg646_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg981_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1038_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg531_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No14_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg626_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No484_out_to_Subtract30_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No485_out_to_Subtract30_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg534_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg963_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg629_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No43_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg775_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No486_out_to_Subtract30_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No487_out_to_Subtract30_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Subtract30_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Subtract30_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Subtract30_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out_to_MUX_Subtract30_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg966_out_to_MUX_Subtract30_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract30_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract30_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg750_out_to_MUX_Subtract30_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg892_out_to_MUX_Subtract30_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Subtract30_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg891_out_to_MUX_Subtract30_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out_to_MUX_Subtract30_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Subtract30_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Subtract30_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out_to_MUX_Subtract30_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Subtract30_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out_to_MUX_Subtract30_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract30_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract30_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Subtract30_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg967_out_to_MUX_Subtract30_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Subtract30_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg966_out_to_MUX_Subtract30_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Subtract30_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No488_out_to_Subtract30_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No489_out_to_Subtract30_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg582_out_to_MUX_Subtract30_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out_to_MUX_Subtract30_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Subtract30_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg991_out_to_MUX_Subtract30_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out_to_MUX_Subtract30_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg969_out_to_MUX_Subtract30_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Subtract30_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract30_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg897_out_to_MUX_Subtract30_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg896_out_to_MUX_Subtract30_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Subtract30_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg895_out_to_MUX_Subtract30_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_Subtract30_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Subtract30_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Subtract30_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No17_out_to_MUX_Subtract30_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out_to_MUX_Subtract30_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg925_out_to_MUX_Subtract30_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract30_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract30_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No45_out_to_MUX_Subtract30_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg970_out_to_MUX_Subtract30_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Subtract30_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg969_out_to_MUX_Subtract30_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No490_out_to_Subtract30_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No491_out_to_Subtract30_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Subtract30_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Subtract30_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Subtract30_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out_to_MUX_Subtract30_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Subtract30_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Subtract30_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Subtract30_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg587_out_to_MUX_Subtract30_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract30_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract30_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Subtract30_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Subtract30_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg994_out_to_MUX_Subtract30_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg972_out_to_MUX_Subtract30_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Subtract30_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_Subtract30_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Subtract30_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Subtract30_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out_to_MUX_Subtract30_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg763_out_to_MUX_Subtract30_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract30_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract30_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Subtract30_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Subtract30_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No492_out_to_Subtract30_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No493_out_to_Subtract30_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Subtract30_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Subtract30_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Subtract30_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out_to_MUX_Subtract30_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Subtract30_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Subtract30_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Subtract30_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Subtract30_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out_to_MUX_Subtract30_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg592_out_to_MUX_Subtract30_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract30_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract30_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Subtract30_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg976_out_to_MUX_Subtract30_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Subtract30_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Subtract30_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Subtract30_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_Subtract30_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out_to_MUX_Subtract30_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Subtract30_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out_to_MUX_Subtract30_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out_to_MUX_Subtract30_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract30_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract30_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No494_out_to_Subtract30_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No495_out_to_Subtract30_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract30_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Subtract30_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Subtract30_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Subtract30_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Subtract30_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out_to_MUX_Subtract30_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out_to_MUX_Subtract30_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out_to_MUX_Subtract30_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Subtract30_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out_to_MUX_Subtract30_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg978_out_to_MUX_Subtract30_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Subtract30_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract30_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Subtract30_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Subtract30_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Subtract30_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Subtract30_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Subtract30_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Subtract30_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Subtract30_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Subtract30_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg644_out_to_MUX_Subtract30_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Subtract30_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract30_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No496_out_to_Subtract32_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No497_out_to_Subtract32_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out_to_MUX_Subtract32_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract32_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract32_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_Subtract32_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Subtract32_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Subtract32_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out_to_MUX_Subtract32_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Subtract32_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Subtract32_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Subtract32_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Subtract32_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out_to_MUX_Subtract32_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out_to_MUX_Subtract32_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract32_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract32_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No42_out_to_MUX_Subtract32_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out_to_MUX_Subtract32_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Subtract32_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out_to_MUX_Subtract32_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Subtract32_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Subtract32_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Subtract32_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Subtract32_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg823_out_to_MUX_Subtract32_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No498_out_to_Subtract32_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No499_out_to_Subtract32_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1043_out_to_MUX_Subtract32_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out_to_MUX_Subtract32_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg676_out_to_MUX_Subtract32_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract32_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract32_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out_to_MUX_Subtract32_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out_to_MUX_Subtract32_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Subtract32_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_Subtract32_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Subtract32_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Subtract32_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg984_out_to_MUX_Subtract32_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1046_out_to_MUX_Subtract32_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out_to_MUX_Subtract32_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out_to_MUX_Subtract32_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract32_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract32_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Subtract32_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg964_out_to_MUX_Subtract32_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Subtract32_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg963_out_to_MUX_Subtract32_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Subtract32_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Subtract32_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out_to_MUX_Subtract32_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No500_out_to_Subtract32_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No501_out_to_Subtract32_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out_to_MUX_Subtract32_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Subtract32_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1013_out_to_MUX_Subtract32_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Subtract32_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg682_out_to_MUX_Subtract32_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract32_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract32_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Subtract32_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out_to_MUX_Subtract32_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out_to_MUX_Subtract32_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Subtract32_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Subtract32_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Subtract32_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg751_out_to_MUX_Subtract32_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1016_out_to_MUX_Subtract32_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out_to_MUX_Subtract32_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out_to_MUX_Subtract32_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract32_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract32_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Subtract32_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Subtract32_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg987_out_to_MUX_Subtract32_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Subtract32_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Subtract32_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No502_out_to_Subtract32_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No503_out_to_Subtract32_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Subtract32_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Subtract32_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Subtract32_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Subtract32_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out_to_MUX_Subtract32_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out_to_MUX_Subtract32_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract32_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract32_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out_to_MUX_Subtract32_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg880_out_to_MUX_Subtract32_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out_to_MUX_Subtract32_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Subtract32_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Subtract32_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Subtract32_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg756_out_to_MUX_Subtract32_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out_to_MUX_Subtract32_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Subtract32_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Subtract32_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract32_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract32_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out_to_MUX_Subtract32_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out_to_MUX_Subtract32_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg991_out_to_MUX_Subtract32_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Subtract32_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No504_out_to_Subtract32_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No505_out_to_Subtract32_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Subtract32_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out_to_MUX_Subtract32_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Subtract32_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Subtract32_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out_to_MUX_Subtract32_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Subtract32_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Subtract32_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1029_out_to_MUX_Subtract32_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out_to_MUX_Subtract32_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Subtract32_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract32_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract32_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Subtract32_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Subtract32_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_Subtract32_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg975_out_to_MUX_Subtract32_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out_to_MUX_Subtract32_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Subtract32_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Subtract32_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1065_out_to_MUX_Subtract32_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Subtract32_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Subtract32_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract32_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract32_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No506_out_to_Subtract32_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No507_out_to_Subtract32_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract32_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Subtract32_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Subtract32_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Subtract32_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Subtract32_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Subtract32_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Subtract32_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Subtract32_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1034_out_to_MUX_Subtract32_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out_to_MUX_Subtract32_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg703_out_to_MUX_Subtract32_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract32_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract32_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No48_out_to_MUX_Subtract32_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg979_out_to_MUX_Subtract32_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out_to_MUX_Subtract32_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out_to_MUX_Subtract32_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Subtract32_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Subtract32_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Subtract32_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No20_out_to_MUX_Subtract32_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out_to_MUX_Subtract32_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out_to_MUX_Subtract32_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract32_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No508_out_to_Subtract43_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No509_out_to_Subtract43_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out_to_MUX_Subtract43_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract43_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract43_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Subtract43_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out_to_MUX_Subtract43_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Subtract43_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Subtract43_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Subtract43_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Subtract43_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1004_out_to_MUX_Subtract43_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1071_out_to_MUX_Subtract43_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Subtract43_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Subtract43_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract43_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract43_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Subtract43_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg961_out_to_MUX_Subtract43_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Subtract43_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg960_out_to_MUX_Subtract43_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg666_out_to_MUX_Subtract43_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Subtract43_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Subtract43_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1074_out_to_MUX_Subtract43_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg960_out_to_MUX_Subtract43_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No510_out_to_Subtract44_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No511_out_to_Subtract44_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract44_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out_to_MUX_Subtract44_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg477_out_to_MUX_Subtract44_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Subtract44_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Subtract44_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out_to_MUX_Subtract44_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg702_out_to_MUX_Subtract44_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1001_out_to_MUX_Subtract44_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Subtract44_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg958_out_to_MUX_Subtract44_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out_to_MUX_Subtract44_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract44_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract44_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out_to_MUX_Subtract44_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out_to_MUX_Subtract44_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Subtract44_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg978_out_to_MUX_Subtract44_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Subtract44_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Subtract44_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg601_out_to_MUX_Subtract44_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out_to_MUX_Subtract44_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg978_out_to_MUX_Subtract44_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out_to_MUX_Subtract44_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract44_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No512_out_to_Subtract49_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No513_out_to_Subtract49_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Subtract49_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Subtract49_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Subtract49_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract49_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract49_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Subtract49_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out_to_MUX_Subtract49_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Subtract49_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Subtract49_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Subtract49_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Subtract49_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Subtract49_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out_to_MUX_Subtract49_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg963_out_to_MUX_Subtract49_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Subtract49_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract49_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract49_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Subtract49_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Subtract49_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg985_out_to_MUX_Subtract49_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Subtract49_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Subtract49_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg984_out_to_MUX_Subtract49_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Subtract49_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No514_out_to_Subtract116_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No515_out_to_Subtract116_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract116_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Subtract116_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg874_out_to_MUX_Subtract116_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg703_out_to_MUX_Subtract116_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg360_out_to_MUX_Subtract116_6_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Subtract116_6_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Subtract116_6_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Subtract116_6_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1067_out_to_MUX_Subtract116_6_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Subtract116_6_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg873_out_to_MUX_Subtract116_6_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract116_6_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract116_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out_to_MUX_Subtract116_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out_to_MUX_Subtract116_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1002_out_to_MUX_Subtract116_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Subtract116_6_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Subtract116_6_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Subtract116_6_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out_to_MUX_Subtract116_6_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1080_out_to_MUX_Subtract116_6_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Subtract116_6_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg875_out_to_MUX_Subtract116_6_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract116_6_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No516_out_to_Subtract58_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No517_out_to_Subtract58_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out_to_MUX_Subtract58_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract58_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract58_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Subtract58_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Subtract58_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out_to_MUX_Subtract58_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Subtract58_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Subtract58_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Subtract58_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Subtract58_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Subtract58_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out_to_MUX_Subtract58_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out_to_MUX_Subtract58_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract58_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract58_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Subtract58_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Subtract58_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg982_out_to_MUX_Subtract58_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Subtract58_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Subtract58_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1004_out_to_MUX_Subtract58_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Subtract58_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_Subtract58_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Subtract58_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No518_out_to_Subtract125_6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No519_out_to_Subtract125_6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Subtract125_6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out_to_MUX_Subtract125_6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Subtract125_6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out_to_MUX_Subtract125_6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract125_6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Subtract125_6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1033_out_to_MUX_Subtract125_6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Subtract125_6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   ModCount121_instance: ModuloCounter_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Counter_out => ModCount121_out);
x0_re_0_IEEE <= x0_re_0;
   x0_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x0_re_0_out,
                 X => x0_re_0_IEEE);
x0_im_0_IEEE <= x0_im_0;
   x0_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x0_im_0_out,
                 X => x0_im_0_IEEE);
x1_re_0_IEEE <= x1_re_0;
   x1_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x1_re_0_out,
                 X => x1_re_0_IEEE);
x1_im_0_IEEE <= x1_im_0;
   x1_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x1_im_0_out,
                 X => x1_im_0_IEEE);
x2_re_0_IEEE <= x2_re_0;
   x2_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x2_re_0_out,
                 X => x2_re_0_IEEE);
x2_im_0_IEEE <= x2_im_0;
   x2_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x2_im_0_out,
                 X => x2_im_0_IEEE);
x3_re_0_IEEE <= x3_re_0;
   x3_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x3_re_0_out,
                 X => x3_re_0_IEEE);
x3_im_0_IEEE <= x3_im_0;
   x3_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x3_im_0_out,
                 X => x3_im_0_IEEE);
x4_re_0_IEEE <= x4_re_0;
   x4_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x4_re_0_out,
                 X => x4_re_0_IEEE);
x4_im_0_IEEE <= x4_im_0;
   x4_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x4_im_0_out,
                 X => x4_im_0_IEEE);
x5_re_0_IEEE <= x5_re_0;
   x5_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x5_re_0_out,
                 X => x5_re_0_IEEE);
x5_im_0_IEEE <= x5_im_0;
   x5_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x5_im_0_out,
                 X => x5_im_0_IEEE);
x6_re_0_IEEE <= x6_re_0;
   x6_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x6_re_0_out,
                 X => x6_re_0_IEEE);
x6_im_0_IEEE <= x6_im_0;
   x6_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x6_im_0_out,
                 X => x6_im_0_IEEE);
x7_re_0_IEEE <= x7_re_0;
   x7_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x7_re_0_out,
                 X => x7_re_0_IEEE);
x7_im_0_IEEE <= x7_im_0;
   x7_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x7_im_0_out,
                 X => x7_im_0_IEEE);
x8_re_0_IEEE <= x8_re_0;
   x8_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x8_re_0_out,
                 X => x8_re_0_IEEE);
x8_im_0_IEEE <= x8_im_0;
   x8_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x8_im_0_out,
                 X => x8_im_0_IEEE);
x9_re_0_IEEE <= x9_re_0;
   x9_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x9_re_0_out,
                 X => x9_re_0_IEEE);
x9_im_0_IEEE <= x9_im_0;
   x9_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x9_im_0_out,
                 X => x9_im_0_IEEE);
x10_re_0_IEEE <= x10_re_0;
   x10_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x10_re_0_out,
                 X => x10_re_0_IEEE);
x10_im_0_IEEE <= x10_im_0;
   x10_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x10_im_0_out,
                 X => x10_im_0_IEEE);
x11_re_0_IEEE <= x11_re_0;
   x11_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x11_re_0_out,
                 X => x11_re_0_IEEE);
x11_im_0_IEEE <= x11_im_0;
   x11_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x11_im_0_out,
                 X => x11_im_0_IEEE);
x12_re_0_IEEE <= x12_re_0;
   x12_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x12_re_0_out,
                 X => x12_re_0_IEEE);
x12_im_0_IEEE <= x12_im_0;
   x12_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x12_im_0_out,
                 X => x12_im_0_IEEE);
x13_re_0_IEEE <= x13_re_0;
   x13_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x13_re_0_out,
                 X => x13_re_0_IEEE);
x13_im_0_IEEE <= x13_im_0;
   x13_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x13_im_0_out,
                 X => x13_im_0_IEEE);
x14_re_0_IEEE <= x14_re_0;
   x14_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x14_re_0_out,
                 X => x14_re_0_IEEE);
x14_im_0_IEEE <= x14_im_0;
   x14_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x14_im_0_out,
                 X => x14_im_0_IEEE);
x15_re_0_IEEE <= x15_re_0;
   x15_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x15_re_0_out,
                 X => x15_re_0_IEEE);
x15_im_0_IEEE <= x15_im_0;
   x15_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x15_im_0_out,
                 X => x15_im_0_IEEE);
   y0_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y0_re_0_IEEE,
                 X => Delay1No_out);
y0_re_0 <= y0_re_0_IEEE;

SharedReg65_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg65_out;
SharedReg69_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg69_out;
SharedReg105_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg105_out;
SharedReg77_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg77_out;
SharedReg81_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg81_out;
SharedReg118_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg118_out;
SharedReg91_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg91_out;
   MUX_y0_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg65_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg69_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg105_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg77_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg81_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg118_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg91_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y0_re_0_0_LUT_out,
                 oMux => MUX_y0_re_0_0_out);

   Delay1No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y0_re_0_0_out,
                 Y => Delay1No_out);
   y0_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y0_im_0_IEEE,
                 X => Delay1No1_out);
y0_im_0 <= y0_im_0_IEEE;

SharedReg95_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg95_out;
SharedReg100_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg100_out;
SharedReg134_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg134_out;
SharedReg110_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg110_out;
SharedReg114_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg114_out;
SharedReg150_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg150_out;
SharedReg123_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg123_out;
   MUX_y0_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg95_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg100_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg134_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg110_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg114_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg150_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg123_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y0_im_0_0_LUT_out,
                 oMux => MUX_y0_im_0_0_out);

   Delay1No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y0_im_0_0_out,
                 Y => Delay1No1_out);
   y1_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y1_re_0_IEEE,
                 X => Delay1No2_out);
y1_re_0 <= y1_re_0_IEEE;

SharedReg202_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg202_out;
SharedReg130_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg130_out;
SharedReg239_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg239_out;
SharedReg139_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg139_out;
SharedReg206_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg206_out;
SharedReg286_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg286_out;
SharedReg187_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg187_out;
   MUX_y1_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg202_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg239_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg139_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg206_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg286_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg187_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y1_re_0_0_LUT_out,
                 oMux => MUX_y1_re_0_0_out);

   Delay1No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y1_re_0_0_out,
                 Y => Delay1No2_out);
   y1_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y1_im_0_IEEE,
                 X => Delay1No3_out);
y1_im_0 <= y1_im_0_IEEE;

SharedReg249_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg249_out;
SharedReg234_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg234_out;
SharedReg260_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg260_out;
SharedReg244_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg244_out;
SharedReg272_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg272_out;
SharedReg290_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg290_out;
SharedReg218_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg218_out;
   MUX_y1_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg249_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg234_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg260_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg244_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg272_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg290_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg218_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y1_im_0_0_LUT_out,
                 oMux => MUX_y1_im_0_0_out);

   Delay1No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y1_im_0_0_out,
                 Y => Delay1No3_out);
   y2_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y2_re_0_IEEE,
                 X => Delay1No4_out);
y2_re_0 <= y2_re_0_IEEE;

SharedReg65_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg65_out;
SharedReg38_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg38_out;
SharedReg41_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg41_out;
SharedReg198_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg198_out;
SharedReg48_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg48_out;
SharedReg118_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg118_out;
SharedReg91_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg91_out;
   MUX_y2_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg65_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg38_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg41_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg198_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg48_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg118_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg91_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y2_re_0_0_LUT_out,
                 oMux => MUX_y2_re_0_0_out);

   Delay1No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y2_re_0_0_out,
                 Y => Delay1No4_out);
   y2_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y2_im_0_IEEE,
                 X => Delay1No5_out);
y2_im_0 <= y2_im_0_IEEE;

SharedReg95_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg95_out;
SharedReg69_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg69_out;
SharedReg73_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg73_out;
SharedReg44_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg44_out;
SharedReg81_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg81_out;
SharedReg150_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg150_out;
SharedReg123_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg123_out;
   MUX_y2_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg95_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg69_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg73_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg44_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg81_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg150_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg123_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y2_im_0_0_LUT_out,
                 oMux => MUX_y2_im_0_0_out);

   Delay1No5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y2_im_0_0_out,
                 Y => Delay1No5_out);
   y3_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y3_re_0_IEEE,
                 X => Delay1No6_out);
y3_re_0 <= y3_re_0_IEEE;

SharedReg363_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg363_out;
SharedReg372_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg372_out;
SharedReg170_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg170_out;
SharedReg191_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg191_out;
SharedReg52_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg52_out;
SharedReg60_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg60_out;
SharedReg381_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg381_out;
   MUX_y3_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg363_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg372_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg170_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg191_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg52_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg60_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg381_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y3_re_0_0_LUT_out,
                 oMux => MUX_y3_re_0_0_out);

   Delay1No6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y3_re_0_0_out,
                 Y => Delay1No6_out);
   y3_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y3_im_0_IEEE,
                 X => Delay1No7_out);
y3_im_0 <= y3_im_0_IEEE;

SharedReg202_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg202_out;
SharedReg130_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg130_out;
SharedReg239_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg239_out;
SharedReg244_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg244_out;
SharedReg206_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg206_out;
SharedReg212_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg212_out;
SharedReg218_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg218_out;
   MUX_y3_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg202_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg239_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg244_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg206_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg212_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg218_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y3_im_0_0_LUT_out,
                 oMux => MUX_y3_im_0_0_out);

   Delay1No7_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y3_im_0_0_out,
                 Y => Delay1No7_out);
   y4_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y4_re_0_IEEE,
                 X => Delay1No8_out);
y4_re_0 <= y4_re_0_IEEE;

SharedReg127_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg127_out;
SharedReg130_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg130_out;
SharedReg239_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg239_out;
SharedReg139_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg139_out;
SharedReg145_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg145_out;
SharedReg182_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg182_out;
SharedReg153_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg153_out;
   MUX_y4_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg127_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg239_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg139_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg145_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg182_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg153_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y4_re_0_0_LUT_out,
                 oMux => MUX_y4_re_0_0_out);

   Delay1No8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y4_re_0_0_out,
                 Y => Delay1No8_out);
   y4_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y4_im_0_IEEE,
                 X => Delay1No9_out);
y4_im_0 <= y4_im_0_IEEE;

SharedReg202_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg202_out;
SharedReg234_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg234_out;
SharedReg260_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg260_out;
SharedReg244_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg244_out;
SharedReg206_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg206_out;
SharedReg212_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg212_out;
SharedReg187_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg187_out;
   MUX_y4_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg202_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg234_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg260_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg244_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg206_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg212_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg187_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y4_im_0_0_LUT_out,
                 oMux => MUX_y4_im_0_0_out);

   Delay1No9_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y4_im_0_0_out,
                 Y => Delay1No9_out);
   y5_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y5_re_0_IEEE,
                 X => Delay1No10_out);
y5_re_0 <= y5_re_0_IEEE;

SharedReg297_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg297_out;
SharedReg254_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg254_out;
SharedReg302_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg302_out;
SharedReg266_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg266_out;
SharedReg308_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg308_out;
SharedReg313_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg313_out;
SharedReg320_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg320_out;
   MUX_y5_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg297_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg254_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg302_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg266_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg308_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg313_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg320_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y5_re_0_0_LUT_out,
                 oMux => MUX_y5_re_0_0_out);

   Delay1No10_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y5_re_0_0_out,
                 Y => Delay1No10_out);
   y5_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y5_im_0_IEEE,
                 X => Delay1No11_out);
y5_im_0 <= y5_im_0_IEEE;

SharedReg326_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg326_out;
SharedReg335_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg335_out;
SharedReg342_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg342_out;
SharedReg350_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg350_out;
SharedReg278_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg278_out;
SharedReg224_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg224_out;
SharedReg355_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg355_out;
   MUX_y5_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg326_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg335_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg342_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg350_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg278_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg224_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg355_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y5_im_0_0_LUT_out,
                 oMux => MUX_y5_im_0_0_out);

   Delay1No11_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y5_im_0_0_out,
                 Y => Delay1No11_out);
   y6_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y6_re_0_IEEE,
                 X => Delay1No12_out);
y6_re_0 <= y6_re_0_IEEE;

SharedReg127_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg127_out;
SharedReg100_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg100_out;
SharedReg105_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg105_out;
SharedReg77_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg77_out;
SharedReg114_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg114_out;
SharedReg182_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg182_out;
SharedReg153_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg153_out;
   MUX_y6_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg127_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg100_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg105_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg77_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg114_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg182_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg153_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y6_re_0_0_LUT_out,
                 oMux => MUX_y6_re_0_0_out);

   Delay1No12_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y6_re_0_0_out,
                 Y => Delay1No12_out);
   y6_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y6_im_0_IEEE,
                 X => Delay1No13_out);
y6_im_0 <= y6_im_0_IEEE;

SharedReg110_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg110_out;
SharedReg202_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg202_out;
SharedReg130_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg130_out;
SharedReg134_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg134_out;
SharedReg145_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg145_out;
SharedReg212_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg212_out;
SharedReg187_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg187_out;
   MUX_y6_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg110_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg202_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg130_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg134_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg145_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg212_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg187_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y6_im_0_0_LUT_out,
                 oMux => MUX_y6_im_0_0_out);

   Delay1No13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y6_im_0_0_out,
                 Y => Delay1No13_out);
   y7_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y7_re_0_IEEE,
                 X => Delay1No14_out);
y7_re_0 <= y7_re_0_IEEE;

SharedReg249_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg249_out;
SharedReg234_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg234_out;
SharedReg260_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg260_out;
SharedReg266_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg266_out;
SharedReg272_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg272_out;
SharedReg286_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg286_out;
SharedReg320_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg320_out;
   MUX_y7_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg249_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg234_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg260_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg266_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg272_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg286_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg320_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y7_re_0_0_LUT_out,
                 oMux => MUX_y7_re_0_0_out);

   Delay1No14_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y7_re_0_0_out,
                 Y => Delay1No14_out);
   y7_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y7_im_0_IEEE,
                 X => Delay1No15_out);
y7_im_0 <= y7_im_0_IEEE;

SharedReg297_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg297_out;
SharedReg254_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg254_out;
SharedReg302_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg302_out;
SharedReg350_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg350_out;
SharedReg308_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg308_out;
SharedReg290_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg290_out;
SharedReg355_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg355_out;
   MUX_y7_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg297_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg254_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg302_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg350_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg308_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg290_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg355_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y7_im_0_0_LUT_out,
                 oMux => MUX_y7_im_0_0_out);

   Delay1No15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y7_im_0_0_out,
                 Y => Delay1No15_out);
   y8_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y8_re_0_IEEE,
                 X => Delay1No16_out);
y8_re_0 <= y8_re_0_IEEE;

SharedReg1037_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg1037_out;
SharedReg1042_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg1042_out;
SharedReg1047_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg1047_out;
SharedReg1054_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg1054_out;
SharedReg1022_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg1022_out;
SharedReg1028_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg1028_out;
SharedReg1066_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg1066_out;
   MUX_y8_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1037_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1042_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1047_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1054_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1022_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1028_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1066_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y8_re_0_0_LUT_out,
                 oMux => MUX_y8_re_0_0_out);

   Delay1No16_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y8_re_0_0_out,
                 Y => Delay1No16_out);
   y8_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y8_im_0_IEEE,
                 X => Delay1No17_out);
y8_im_0 <= y8_im_0_IEEE;

SharedReg1070_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg1070_out;
SharedReg1081_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg1081_out;
SharedReg876_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg876_out;
SharedReg790_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg790_out;
SharedReg795_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg795_out;
SharedReg1060_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg1060_out;
SharedReg1075_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg1075_out;
   MUX_y8_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1070_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1081_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg876_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg790_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg795_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1060_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1075_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y8_im_0_0_LUT_out,
                 oMux => MUX_y8_im_0_0_out);

   Delay1No17_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y8_im_0_0_out,
                 Y => Delay1No17_out);
   y9_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y9_re_0_IEEE,
                 X => Delay1No18_out);
y9_re_0 <= y9_re_0_IEEE;

SharedReg1004_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg1004_out;
SharedReg984_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg984_out;
SharedReg986_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg986_out;
SharedReg990_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg990_out;
SharedReg993_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg993_out;
SharedReg1028_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg1028_out;
SharedReg1033_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg1033_out;
   MUX_y9_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1004_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg984_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg986_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg990_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg993_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1028_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1033_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y9_re_0_0_LUT_out,
                 oMux => MUX_y9_re_0_0_out);

   Delay1No18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y9_re_0_0_out,
                 Y => Delay1No18_out);
   y9_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y9_im_0_IEEE,
                 X => Delay1No19_out);
y9_im_0 <= y9_im_0_IEEE;

SharedReg1037_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg1037_out;
SharedReg1007_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg1007_out;
SharedReg1012_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg1012_out;
SharedReg1017_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg1017_out;
SharedReg1022_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg1022_out;
SharedReg1060_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg1060_out;
SharedReg1066_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg1066_out;
   MUX_y9_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1037_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1007_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1012_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1017_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1022_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1060_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1066_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y9_im_0_0_LUT_out,
                 oMux => MUX_y9_im_0_0_out);

   Delay1No19_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y9_im_0_0_out,
                 Y => Delay1No19_out);
   y10_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y10_re_0_IEEE,
                 X => Delay1No20_out);
y10_re_0 <= y10_re_0_IEEE;

SharedReg666_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg666_out;
SharedReg570_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg570_out;
SharedReg445_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg445_out;
SharedReg451_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg451_out;
SharedReg458_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg458_out;
SharedReg589_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg589_out;
SharedReg699_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg699_out;
   MUX_y10_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg666_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg570_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg445_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg451_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg458_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg589_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg699_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y10_re_0_0_LUT_out,
                 oMux => MUX_y10_re_0_0_out);

   Delay1No20_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y10_re_0_0_out,
                 Y => Delay1No20_out);
   y10_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y10_im_0_IEEE,
                 X => Delay1No21_out);
y10_im_0 <= y10_im_0_IEEE;

SharedReg849_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg849_out;
SharedReg672_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg672_out;
SharedReg576_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg576_out;
SharedReg580_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg580_out;
SharedReg584_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg584_out;
SharedReg694_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg694_out;
SharedReg871_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg871_out;
   MUX_y10_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg849_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg672_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg576_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg580_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg584_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg694_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg871_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y10_im_0_0_LUT_out,
                 oMux => MUX_y10_im_0_0_out);

   Delay1No21_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y10_im_0_0_out,
                 Y => Delay1No21_out);
   y11_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y11_re_0_IEEE,
                 X => Delay1No22_out);
y11_re_0 <= y11_re_0_IEEE;

SharedReg1004_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg1004_out;
SharedReg984_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg984_out;
SharedReg986_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg986_out;
SharedReg1017_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg1017_out;
SharedReg993_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg993_out;
SharedReg997_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg997_out;
SharedReg1066_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg1066_out;
   MUX_y11_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1004_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg984_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg986_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1017_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg993_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg997_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1066_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y11_re_0_0_LUT_out,
                 oMux => MUX_y11_re_0_0_out);

   Delay1No22_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y11_re_0_0_out,
                 Y => Delay1No22_out);
   y11_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y11_im_0_IEEE,
                 X => Delay1No23_out);
y11_im_0 <= y11_im_0_IEEE;

SharedReg1037_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg1037_out;
SharedReg1007_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg1007_out;
SharedReg1012_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg1012_out;
SharedReg1054_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg1054_out;
SharedReg1022_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg1022_out;
SharedReg1028_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg1028_out;
SharedReg1075_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg1075_out;
   MUX_y11_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1037_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1007_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1012_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1054_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1022_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1028_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1075_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y11_im_0_0_LUT_out,
                 oMux => MUX_y11_im_0_0_out);

   Delay1No23_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y11_im_0_0_out,
                 Y => Delay1No23_out);
   y12_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y12_re_0_IEEE,
                 X => Delay1No24_out);
y12_re_0 <= y12_re_0_IEEE;

SharedReg783_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg783_out;
SharedReg1094_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg1094_out;
SharedReg753_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg753_out;
SharedReg758_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg758_out;
SharedReg764_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg764_out;
SharedReg770_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg770_out;
SharedReg1088_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg1088_out;
   MUX_y12_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg783_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1094_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg753_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg758_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg764_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg770_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1088_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y12_re_0_0_LUT_out,
                 oMux => MUX_y12_re_0_0_out);

   Delay1No24_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y12_re_0_0_out,
                 Y => Delay1No24_out);
   y12_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y12_im_0_IEEE,
                 X => Delay1No25_out);
y12_im_0 <= y12_im_0_IEEE;

SharedReg981_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg981_out;
SharedReg984_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg984_out;
SharedReg986_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg986_out;
SharedReg990_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg990_out;
SharedReg865_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg865_out;
SharedReg868_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg868_out;
SharedReg1001_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg1001_out;
   MUX_y12_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg981_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg984_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg986_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg990_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg865_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg868_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1001_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y12_im_0_0_LUT_out,
                 oMux => MUX_y12_im_0_0_out);

   Delay1No25_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y12_im_0_0_out,
                 Y => Delay1No25_out);
   y13_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y13_re_0_IEEE,
                 X => Delay1No26_out);
y13_re_0 <= y13_re_0_IEEE;

SharedReg1070_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg1070_out;
SharedReg1042_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg1042_out;
SharedReg1047_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg1047_out;
SharedReg1054_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg1054_out;
SharedReg795_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg795_out;
SharedReg770_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg770_out;
SharedReg1075_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg1075_out;
   MUX_y13_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1070_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1042_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1047_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1054_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg795_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg770_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1075_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y13_re_0_0_LUT_out,
                 oMux => MUX_y13_re_0_0_out);

   Delay1No26_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y13_re_0_0_out,
                 Y => Delay1No26_out);
   y13_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y13_im_0_IEEE,
                 X => Delay1No27_out);
y13_im_0 <= y13_im_0_IEEE;

SharedReg1094_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg1094_out;
SharedReg1081_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg1081_out;
SharedReg876_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg876_out;
SharedReg790_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg790_out;
SharedReg764_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg764_out;
SharedReg473_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg473_out;
SharedReg1088_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg1088_out;
   MUX_y13_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1094_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1081_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg876_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg790_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg764_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg473_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1088_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y13_im_0_0_LUT_out,
                 oMux => MUX_y13_im_0_0_out);

   Delay1No27_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y13_im_0_0_out,
                 Y => Delay1No27_out);
   y14_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y14_re_0_IEEE,
                 X => Delay1No28_out);
y14_re_0 <= y14_re_0_IEEE;

SharedReg981_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg981_out;
SharedReg854_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg854_out;
SharedReg678_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg678_out;
SharedReg683_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg683_out;
SharedReg689_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg689_out;
SharedReg868_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg868_out;
SharedReg1001_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg1001_out;
   MUX_y14_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg981_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg854_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg678_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg683_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg689_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg868_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1001_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y14_re_0_0_LUT_out,
                 oMux => MUX_y14_re_0_0_out);

   Delay1No28_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y14_re_0_0_out,
                 Y => Delay1No28_out);
   y14_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y14_im_0_IEEE,
                 X => Delay1No29_out);
y14_im_0 <= y14_im_0_IEEE;

SharedReg1004_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg1004_out;
SharedReg984_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg984_out;
SharedReg858_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg858_out;
SharedReg861_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg861_out;
SharedReg865_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg865_out;
SharedReg997_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg997_out;
SharedReg1033_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg1033_out;
   MUX_y14_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1004_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg984_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg858_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg861_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg865_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg997_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1033_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y14_im_0_0_LUT_out,
                 oMux => MUX_y14_im_0_0_out);

   Delay1No29_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y14_im_0_0_out,
                 Y => Delay1No29_out);
   y15_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y15_re_0_IEEE,
                 X => Delay1No30_out);
y15_re_0 <= y15_re_0_IEEE;

SharedReg1060_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg1060_out;
SharedReg795_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg795_out;
SharedReg1070_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg1070_out;
SharedReg1042_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg1042_out;
SharedReg1047_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg1047_out;
SharedReg790_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_6_cast <= SharedReg790_out;
SharedReg1088_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_7_cast <= SharedReg1088_out;
   MUX_y15_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1060_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg795_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1070_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1042_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1047_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg790_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1088_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y15_re_0_0_LUT_out,
                 oMux => MUX_y15_re_0_0_out);

   Delay1No30_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y15_re_0_0_out,
                 Y => Delay1No30_out);
   y15_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y15_im_0_IEEE,
                 X => Delay1No31_out);
y15_im_0 <= y15_im_0_IEEE;

SharedReg1094_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg1094_out;
SharedReg1081_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg1081_out;
SharedReg876_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg876_out;
SharedReg758_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg758_out;
SharedReg764_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg764_out;
SharedReg770_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_6_cast <= SharedReg770_out;
SharedReg1101_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_7_cast <= SharedReg1101_out;
   MUX_y15_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_7_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1094_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1081_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg876_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg758_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg764_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg770_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1101_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_7_cast,
                 iSel => MUX_y15_im_0_0_LUT_out,
                 oMux => MUX_y15_im_0_0_out);

   Delay1No31_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y15_im_0_0_out,
                 Y => Delay1No31_out);

Delay1No32_out_to_Add2_0_impl_parent_implementedSystem_port_0_cast <= Delay1No32_out;
Delay1No33_out_to_Add2_0_impl_parent_implementedSystem_port_1_cast <= Delay1No33_out;
   Add2_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_0_impl_out,
                 X => Delay1No32_out_to_Add2_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No33_out_to_Add2_0_impl_parent_implementedSystem_port_1_cast);

Delay15No_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_1_cast <= Delay15No_out;
SharedReg_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg_out;
SharedReg12_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg12_out;
SharedReg567_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg567_out;
SharedReg435_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg435_out;
SharedReg1004_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1004_out;
SharedReg332_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg332_out;
SharedReg564_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg564_out;
SharedReg99_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg99_out;
SharedReg666_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg666_out;
SharedReg431_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg431_out;
SharedReg395_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg395_out;
   MUX_Add2_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay15No_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg431_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg395_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg12_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg567_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg435_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1004_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg332_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg564_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg99_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg666_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add2_0_impl_0_out);

   Delay1No32_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_0_impl_0_out,
                 Y => Delay1No32_out);

SharedReg368_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg368_out;
SharedReg16_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg16_out;
SharedReg28_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg28_out;
SharedReg432_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg432_out;
SharedReg432_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg432_out;
SharedReg564_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg564_out;
SharedReg203_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg203_out;
SharedReg849_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg849_out;
SharedReg202_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg202_out;
SharedReg982_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg982_out;
SharedReg564_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg564_out;
SharedReg417_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg417_out;
   MUX_Add2_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg368_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg16_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg564_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg417_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg28_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg432_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg432_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg564_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg203_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg849_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg202_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg982_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add2_0_impl_1_out);

   Delay1No33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_0_impl_1_out,
                 Y => Delay1No33_out);

Delay1No34_out_to_Add2_1_impl_parent_implementedSystem_port_0_cast <= Delay1No34_out;
Delay1No35_out_to_Add2_1_impl_parent_implementedSystem_port_1_cast <= Delay1No35_out;
   Add2_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_1_impl_out,
                 X => Delay1No34_out_to_Add2_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No35_out_to_Add2_1_impl_parent_implementedSystem_port_1_cast);

SharedReg70_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg70_out;
SharedReg398_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg398_out;
Delay15No1_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_3_cast <= Delay15No1_out;
SharedReg_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg_out;
SharedReg12_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg12_out;
SharedReg104_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg104_out;
SharedReg677_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg677_out;
SharedReg373_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg373_out;
SharedReg1009_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1009_out;
SharedReg1084_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1084_out;
SharedReg779_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg779_out;
SharedReg438_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg438_out;
   MUX_Add2_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg70_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg398_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg779_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg438_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => Delay15No1_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg12_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg104_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg677_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg373_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1009_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1084_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add2_1_impl_0_out);

   Delay1No34_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_1_impl_0_out,
                 Y => Delay1No34_out);

SharedReg254_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg254_out;
SharedReg419_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg419_out;
SharedReg377_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg377_out;
SharedReg16_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg16_out;
SharedReg28_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg28_out;
SharedReg256_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg256_out;
SharedReg440_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg440_out;
SharedReg335_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg335_out;
SharedReg444_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg444_out;
SharedReg438_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg438_out;
SharedReg1007_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1007_out;
SharedReg571_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg571_out;
   MUX_Add2_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg254_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg419_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1007_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg571_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg377_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg16_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg28_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg256_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg440_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg335_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg444_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg438_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add2_1_impl_1_out);

   Delay1No35_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_1_impl_1_out,
                 Y => Delay1No35_out);

Delay1No36_out_to_Add2_2_impl_parent_implementedSystem_port_0_cast <= Delay1No36_out;
Delay1No37_out_to_Add2_2_impl_parent_implementedSystem_port_1_cast <= Delay1No37_out;
   Add2_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_2_impl_out,
                 X => Delay1No36_out_to_Add2_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No37_out_to_Add2_2_impl_parent_implementedSystem_port_1_cast);

SharedReg749_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg749_out;
SharedReg445_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg445_out;
SharedReg784_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg784_out;
SharedReg15_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg15_out;
SharedReg723_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg723_out;
SharedReg_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg_out;
SharedReg12_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg12_out;
SharedReg109_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg109_out;
SharedReg579_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg579_out;
SharedReg171_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg171_out;
SharedReg1014_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1014_out;
SharedReg879_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg879_out;
   MUX_Add2_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg749_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg445_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1014_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg879_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg784_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg15_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg723_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg12_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg109_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg579_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg171_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add2_2_impl_0_out);

   Delay1No36_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_2_impl_0_out,
                 Y => Delay1No36_out);

SharedReg986_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg986_out;
SharedReg679_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg679_out;
SharedReg746_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg746_out;
SharedReg31_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg31_out;
SharedReg804_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg804_out;
SharedReg16_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg16_out;
SharedReg28_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg28_out;
SharedReg262_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg262_out;
SharedReg748_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg748_out;
SharedReg342_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg342_out;
SharedReg752_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg752_out;
SharedReg746_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg746_out;
   MUX_Add2_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg986_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg679_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg752_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg746_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg746_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg31_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg804_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg16_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg28_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg262_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg748_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg342_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add2_2_impl_1_out);

   Delay1No37_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_2_impl_1_out,
                 Y => Delay1No37_out);

Delay1No38_out_to_Add2_3_impl_parent_implementedSystem_port_0_cast <= Delay1No38_out;
Delay1No39_out_to_Add2_3_impl_parent_implementedSystem_port_1_cast <= Delay1No39_out;
   Add2_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_3_impl_out,
                 X => Delay1No38_out_to_Add2_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No39_out_to_Add2_3_impl_parent_implementedSystem_port_1_cast);

SharedReg178_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg178_out;
SharedReg455_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg455_out;
SharedReg753_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg753_out;
SharedReg877_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg877_out;
SharedReg404_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg404_out;
Delay15No3_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_6_cast <= Delay15No3_out;
SharedReg_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg_out;
SharedReg7_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg7_out;
SharedReg113_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg113_out;
SharedReg422_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg422_out;
SharedReg451_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg451_out;
SharedReg267_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg267_out;
   MUX_Add2_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg178_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg455_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg451_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg267_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg753_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg877_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg404_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay15No3_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg7_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg113_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg422_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add2_3_impl_0_out);

   Delay1No38_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_3_impl_0_out,
                 Y => Delay1No38_out);

SharedReg266_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg266_out;
SharedReg1017_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1017_out;
SharedReg581_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg581_out;
SharedReg753_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg753_out;
SharedReg423_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg423_out;
Delay10No3_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_6_cast <= Delay10No3_out;
SharedReg16_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg16_out;
SharedReg23_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg23_out;
SharedReg267_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg267_out;
SharedReg489_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg489_out;
SharedReg862_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg862_out;
SharedReg271_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg271_out;
   MUX_Add2_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg266_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1017_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg862_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg271_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg581_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg753_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg423_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay10No3_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg16_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg23_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg267_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg489_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add2_3_impl_1_out);

   Delay1No39_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_3_impl_1_out,
                 Y => Delay1No39_out);

Delay1No40_out_to_Add2_4_impl_parent_implementedSystem_port_0_cast <= Delay1No40_out;
Delay1No41_out_to_Add2_4_impl_parent_implementedSystem_port_1_cast <= Delay1No41_out;
   Add2_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_4_impl_out,
                 X => Delay1No40_out_to_Add2_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No41_out_to_Add2_4_impl_parent_implementedSystem_port_1_cast);

SharedReg705_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg705_out;
SharedReg1023_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1023_out;
SharedReg767_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg767_out;
SharedReg148_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg148_out;
SharedReg705_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg705_out;
SharedReg791_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg791_out;
SharedReg15_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg15_out;
Delay15No4_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_8_cast <= Delay15No4_out;
SharedReg_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg_out;
SharedReg7_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg7_out;
SharedReg210_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg210_out;
SharedReg424_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg424_out;
   MUX_Add2_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg705_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1023_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg210_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg424_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg767_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg148_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg705_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg791_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg15_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay15No4_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg7_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add2_4_impl_0_out);

   Delay1No40_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_4_impl_0_out,
                 Y => Delay1No40_out);

SharedReg866_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg866_out;
SharedReg711_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg711_out;
SharedReg758_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg758_out;
SharedReg114_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg114_out;
SharedReg585_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg585_out;
SharedReg758_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg758_out;
SharedReg31_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg31_out;
SharedReg58_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg58_out;
SharedReg16_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg16_out;
SharedReg23_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg23_out;
SharedReg280_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg280_out;
SharedReg492_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg492_out;
   MUX_Add2_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg866_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg711_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg280_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg492_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg758_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg114_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg585_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg758_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg31_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg58_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg16_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg23_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add2_4_impl_1_out);

   Delay1No41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_4_impl_1_out,
                 Y => Delay1No41_out);

Delay1No42_out_to_Add2_5_impl_parent_implementedSystem_port_0_cast <= Delay1No42_out;
Delay1No43_out_to_Add2_5_impl_parent_implementedSystem_port_1_cast <= Delay1No43_out;
   Add2_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_5_impl_out,
                 X => Delay1No42_out_to_Add2_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No43_out_to_Add2_5_impl_parent_implementedSystem_port_1_cast);

SharedReg122_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg122_out;
SharedReg768_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg768_out;
SharedReg997_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg997_out;
SharedReg928_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg928_out;
SharedReg865_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg865_out;
SharedReg638_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg638_out;
SharedReg927_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg927_out;
SharedReg930_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg930_out;
SharedReg13_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg13_out;
SharedReg735_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg735_out;
SharedReg_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg_out;
SharedReg12_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg12_out;
   MUX_Add2_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg122_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg768_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg12_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg997_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg928_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg865_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg638_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg927_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg930_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg13_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg735_out_to_MUX_Add2_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add2_5_impl_0_out);

   Delay1No42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_5_impl_0_out,
                 Y => Delay1No42_out);

SharedReg292_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg292_out;
SharedReg466_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg466_out;
SharedReg464_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg464_out;
SharedReg952_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg952_out;
SharedReg996_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg996_out;
SharedReg409_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg409_out;
SharedReg900_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg900_out;
Delay4No263_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_8_cast <= Delay4No263_out;
SharedReg29_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg29_out;
SharedReg813_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg813_out;
SharedReg16_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg16_out;
SharedReg28_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg28_out;
   MUX_Add2_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg292_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg466_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg16_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg28_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg464_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg952_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg996_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg409_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg900_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay4No263_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg29_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg813_out_to_MUX_Add2_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add2_5_impl_1_out);

   Delay1No43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_5_impl_1_out,
                 Y => Delay1No43_out);

Delay1No44_out_to_Add2_6_impl_parent_implementedSystem_port_0_cast <= Delay1No44_out;
Delay1No45_out_to_Add2_6_impl_parent_implementedSystem_port_1_cast <= Delay1No45_out;
   Add2_6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_6_impl_out,
                 X => Delay1No44_out_to_Add2_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No45_out_to_Add2_6_impl_parent_implementedSystem_port_1_cast);

SharedReg7_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg7_out;
SharedReg600_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg600_out;
SharedReg874_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg874_out;
SharedReg1033_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1033_out;
SharedReg360_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg360_out;
SharedReg473_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg473_out;
SharedReg997_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg997_out;
SharedReg595_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg595_out;
SharedReg976_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg976_out;
SharedReg413_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg413_out;
Delay15No6_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_11_cast <= Delay15No6_out;
SharedReg_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg_out;
   MUX_Add2_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg7_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg600_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay15No6_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg874_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1033_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg360_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg473_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg997_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg595_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg976_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg413_out_to_MUX_Add2_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add2_6_impl_0_out);

   Delay1No44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_6_impl_0_out,
                 Y => Delay1No44_out);

SharedReg23_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg23_out;
SharedReg597_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg597_out;
SharedReg701_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg701_out;
SharedReg595_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg595_out;
SharedReg189_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg189_out;
SharedReg699_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg699_out;
SharedReg1032_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1032_out;
SharedReg1002_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1002_out;
SharedReg954_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg954_out;
SharedReg429_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg429_out;
SharedReg393_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg393_out;
SharedReg16_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg16_out;
   MUX_Add2_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg23_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg597_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg393_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg16_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg701_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg595_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg189_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg699_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1032_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1002_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg954_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg429_out_to_MUX_Add2_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add2_6_impl_1_out);

   Delay1No45_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_6_impl_1_out,
                 Y => Delay1No45_out);

Delay1No46_out_to_Add11_0_impl_parent_implementedSystem_port_0_cast <= Delay1No46_out;
Delay1No47_out_to_Add11_0_impl_parent_implementedSystem_port_1_cast <= Delay1No47_out;
   Add11_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_0_impl_out,
                 X => Delay1No46_out_to_Add11_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No47_out_to_Add11_0_impl_parent_implementedSystem_port_1_cast);

SharedReg669_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg669_out;
SharedReg1_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1_out;
SharedReg7_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg7_out;
SharedReg129_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg129_out;
SharedReg853_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg853_out;
SharedReg327_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg327_out;
SharedReg1006_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1006_out;
SharedReg1073_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1073_out;
SharedReg434_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg434_out;
SharedReg564_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg564_out;
SharedReg96_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg96_out;
SharedReg501_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg501_out;
   MUX_Add11_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg669_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg96_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg501_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg7_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg129_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg853_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg327_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1006_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1073_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg434_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg564_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add11_0_impl_0_out);

   Delay1No46_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_0_impl_0_out,
                 Y => Delay1No46_out);

SharedReg437_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg437_out;
SharedReg17_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg17_out;
SharedReg23_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg23_out;
SharedReg298_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg298_out;
SharedReg566_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg566_out;
SharedReg297_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg297_out;
SharedReg569_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg569_out;
SharedReg430_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg430_out;
SharedReg1037_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1037_out;
SharedReg667_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg667_out;
SharedReg297_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg297_out;
SharedReg529_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg529_out;
   MUX_Add11_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg437_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg17_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg297_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg529_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg23_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg298_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg566_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg297_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg569_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg430_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1037_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg667_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add11_0_impl_1_out);

   Delay1No47_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_0_impl_1_out,
                 Y => Delay1No47_out);

Delay1No48_out_to_Add11_1_impl_parent_implementedSystem_port_0_cast <= Delay1No48_out;
Delay1No49_out_to_Add11_1_impl_parent_implementedSystem_port_1_cast <= Delay1No49_out;
   Add11_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_1_impl_out,
                 X => Delay1No48_out_to_Add11_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No49_out_to_Add11_1_impl_parent_implementedSystem_port_1_cast);

SharedReg673_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg673_out;
SharedReg505_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg505_out;
SharedReg676_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg676_out;
SharedReg1_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1_out;
SharedReg7_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg7_out;
SharedReg257_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg257_out;
SharedReg418_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg418_out;
SharedReg438_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg438_out;
SharedReg256_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg256_out;
SharedReg166_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg166_out;
SharedReg338_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg338_out;
SharedReg100_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg100_out;
   MUX_Add11_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg673_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg505_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg338_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg100_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg676_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg7_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg257_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg418_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg438_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg256_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg166_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add11_1_impl_0_out);

   Delay1No48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_1_impl_0_out,
                 Y => Delay1No48_out);

SharedReg672_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg672_out;
SharedReg532_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg532_out;
SharedReg782_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg782_out;
SharedReg17_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg17_out;
SharedReg23_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg23_out;
SharedReg337_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg337_out;
SharedReg483_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg483_out;
SharedReg855_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg855_out;
SharedReg341_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg341_out;
SharedReg335_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg335_out;
SharedReg372_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg372_out;
SharedReg235_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg235_out;
   MUX_Add11_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg672_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg532_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg372_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg235_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg782_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg17_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg23_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg337_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg483_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg855_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg341_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg335_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add11_1_impl_1_out);

   Delay1No49_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_1_impl_1_out,
                 Y => Delay1No49_out);

Delay1No50_out_to_Add11_2_impl_parent_implementedSystem_port_0_cast <= Delay1No50_out;
Delay1No51_out_to_Add11_2_impl_parent_implementedSystem_port_1_cast <= Delay1No51_out;
   Add11_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_2_impl_out,
                 X => Delay1No50_out_to_Add11_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No51_out_to_Add11_2_impl_parent_implementedSystem_port_1_cast);

SharedReg346_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg346_out;
SharedReg746_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg746_out;
SharedReg74_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg74_out;
SharedReg401_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg401_out;
Delay15No2_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_5_cast <= Delay15No2_out;
SharedReg1_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1_out;
SharedReg7_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg7_out;
SharedReg263_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg263_out;
SharedReg420_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg420_out;
SharedReg445_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg445_out;
SharedReg304_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg304_out;
SharedReg200_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg200_out;
   MUX_Add11_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg346_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg746_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg304_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg200_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg74_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg401_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay15No2_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg7_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg263_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg420_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg445_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add11_2_impl_0_out);

   Delay1No50_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_2_impl_0_out,
                 Y => Delay1No50_out);

SharedReg342_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg342_out;
SharedReg446_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg446_out;
SharedReg260_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg260_out;
SharedReg421_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg421_out;
Delay10No2_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_5_cast <= Delay10No2_out;
SharedReg17_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg17_out;
SharedReg23_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg23_out;
SharedReg304_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg304_out;
SharedReg486_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg486_out;
SharedReg859_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg859_out;
SharedReg307_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg307_out;
SharedReg302_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg302_out;
   MUX_Add11_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg342_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg446_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg307_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg302_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg260_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg421_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay10No2_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg17_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg23_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg304_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg486_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg859_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add11_2_impl_1_out);

   Delay1No51_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_2_impl_1_out,
                 Y => Delay1No51_out);

Delay1No52_out_to_Add11_3_impl_parent_implementedSystem_port_0_cast <= Delay1No52_out;
Delay1No53_out_to_Add11_3_impl_parent_implementedSystem_port_1_cast <= Delay1No53_out;
   Add11_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_3_impl_out,
                 X => Delay1No52_out_to_Add11_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No53_out_to_Add11_3_impl_parent_implementedSystem_port_1_cast);

SharedReg47_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg47_out;
SharedReg194_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg194_out;
SharedReg77_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg77_out;
SharedReg45_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg45_out;
SharedReg513_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg513_out;
SharedReg687_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg687_out;
SharedReg1_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1_out;
SharedReg8_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg8_out;
SharedReg268_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg268_out;
SharedReg556_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg556_out;
SharedReg266_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg266_out;
SharedReg1055_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1055_out;
   MUX_Add11_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg47_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg194_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg266_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1055_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg77_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg45_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg513_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg687_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg8_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg268_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg556_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add11_3_impl_0_out);

   Delay1No52_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_3_impl_0_out,
                 Y => Delay1No52_out);

SharedReg191_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg191_out;
SharedReg191_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg191_out;
SharedReg245_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg245_out;
SharedReg244_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg244_out;
SharedReg538_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg538_out;
SharedReg882_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg882_out;
SharedReg17_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg17_out;
SharedReg24_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg24_out;
SharedReg352_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg352_out;
SharedReg612_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg612_out;
SharedReg140_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg140_out;
SharedReg457_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg457_out;
   MUX_Add11_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg191_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg191_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg140_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg457_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg245_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg244_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg538_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg882_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg17_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg24_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg352_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg612_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add11_3_impl_1_out);

   Delay1No53_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_3_impl_1_out,
                 Y => Delay1No53_out);

Delay1No54_out_to_Add11_4_impl_parent_implementedSystem_port_0_cast <= Delay1No54_out;
Delay1No55_out_to_Add11_4_impl_parent_implementedSystem_port_1_cast <= Delay1No55_out;
   Add11_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_4_impl_out,
                 X => Delay1No54_out_to_Add11_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No55_out_to_Add11_4_impl_parent_implementedSystem_port_1_cast);

SharedReg272_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg272_out;
SharedReg310_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg310_out;
SharedReg89_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg89_out;
SharedReg708_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg708_out;
SharedReg758_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg758_out;
SharedReg49_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg49_out;
SharedReg407_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg407_out;
SharedReg587_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg587_out;
SharedReg1_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1_out;
SharedReg8_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg8_out;
SharedReg425_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg425_out;
SharedReg558_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg558_out;
   MUX_Add11_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg272_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg310_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg425_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg558_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg89_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg708_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg758_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg49_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg407_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg587_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg8_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add11_4_impl_0_out);

   Delay1No54_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_4_impl_0_out,
                 Y => Delay1No54_out);

SharedReg207_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg207_out;
SharedReg312_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg312_out;
SharedReg272_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg272_out;
SharedReg865_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg865_out;
SharedReg706_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg706_out;
SharedReg206_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg206_out;
SharedReg425_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg425_out;
SharedReg763_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg763_out;
SharedReg17_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg17_out;
SharedReg24_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg24_out;
SharedReg493_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg493_out;
SharedReg615_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg615_out;
   MUX_Add11_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg207_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg312_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg493_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg615_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg272_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg865_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg706_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg206_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg425_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg763_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg17_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg24_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add11_4_impl_1_out);

   Delay1No55_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_4_impl_1_out,
                 Y => Delay1No55_out);

Delay1No56_out_to_Add11_5_impl_parent_implementedSystem_port_0_cast <= Delay1No56_out;
Delay1No57_out_to_Add11_5_impl_parent_implementedSystem_port_1_cast <= Delay1No57_out;
   Add11_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_5_impl_out,
                 X => Delay1No56_out_to_Add11_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No57_out_to_Add11_5_impl_parent_implementedSystem_port_1_cast);

SharedReg216_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg216_out;
SharedReg470_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg470_out;
SharedReg225_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg225_out;
SharedReg294_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg294_out;
SharedReg712_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg712_out;
SharedReg185_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg185_out;
SharedReg973_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg973_out;
SharedReg765_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg765_out;
SharedReg15_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg15_out;
Delay15No5_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_10_cast <= Delay15No5_out;
SharedReg1_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1_out;
SharedReg7_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg7_out;
   MUX_Add11_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg216_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg470_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg7_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg225_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg294_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg712_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg185_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg973_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg765_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg15_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay15No5_out_to_MUX_Add11_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add11_5_impl_0_out);

   Delay1No56_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_5_impl_0_out,
                 Y => Delay1No56_out);

SharedReg315_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg315_out;
SharedReg467_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg467_out;
SharedReg290_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg290_out;
SharedReg288_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg288_out;
SharedReg589_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg589_out;
SharedReg150_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg150_out;
SharedReg951_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg951_out;
SharedReg712_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg712_out;
SharedReg31_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg31_out;
SharedReg230_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg230_out;
SharedReg17_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg17_out;
SharedReg23_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg23_out;
   MUX_Add11_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg315_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg467_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg17_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg23_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg290_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg288_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg589_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg150_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg951_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg712_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg31_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg230_out_to_MUX_Add11_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add11_5_impl_1_out);

   Delay1No57_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_5_impl_1_out,
                 Y => Delay1No57_out);

Delay1No58_out_to_Add11_6_impl_parent_implementedSystem_port_0_cast <= Delay1No58_out;
Delay1No59_out_to_Add11_6_impl_parent_implementedSystem_port_1_cast <= Delay1No59_out;
   Add11_6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_6_impl_out,
                 X => Delay1No58_out_to_Add11_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No59_out_to_Add11_6_impl_parent_implementedSystem_port_1_cast);

SharedReg8_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg8_out;
SharedReg157_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg157_out;
SharedReg428_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg428_out;
SharedReg356_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg356_out;
SharedReg1035_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1035_out;
SharedReg1078_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1078_out;
SharedReg126_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg126_out;
SharedReg473_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg473_out;
SharedReg771_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg771_out;
SharedReg525_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg525_out;
SharedReg703_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg703_out;
SharedReg1_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1_out;
   MUX_Add11_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg8_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg157_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg703_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg428_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg356_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1035_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1078_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg126_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg473_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg771_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg525_out_to_MUX_Add11_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add11_6_impl_0_out);

   Delay1No58_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_6_impl_0_out,
                 Y => Delay1No58_out);

SharedReg24_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg24_out;
SharedReg357_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg357_out;
SharedReg498_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg498_out;
SharedReg320_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg320_out;
SharedReg602_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg602_out;
SharedReg770_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg770_out;
SharedReg187_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg187_out;
SharedReg700_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg700_out;
SharedReg595_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg595_out;
SharedReg547_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg547_out;
SharedReg479_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg479_out;
SharedReg17_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg17_out;
   MUX_Add11_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg24_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg357_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg479_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg17_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg498_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg320_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg602_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg770_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg187_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg700_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg595_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg547_out_to_MUX_Add11_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add11_6_impl_1_out);

   Delay1No59_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_6_impl_1_out,
                 Y => Delay1No59_out);

Delay1No60_out_to_Add3_0_impl_parent_implementedSystem_port_0_cast <= Delay1No60_out;
Delay1No61_out_to_Add3_0_impl_parent_implementedSystem_port_1_cast <= Delay1No61_out;
   Add3_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add3_0_impl_out,
                 X => Delay1No60_out_to_Add3_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No61_out_to_Add3_0_impl_parent_implementedSystem_port_1_cast);

SharedReg331_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg331_out;
SharedReg2_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg2_out;
SharedReg8_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg8_out;
SharedReg299_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg299_out;
SharedReg416_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg416_out;
SharedReg430_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg430_out;
SharedReg251_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg251_out;
SharedReg365_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg365_out;
SharedReg330_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg330_out;
SharedReg127_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg127_out;
SharedReg850_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg850_out;
SharedReg481_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg481_out;
   MUX_Add3_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg331_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg2_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg850_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg481_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg8_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg299_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg416_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg430_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg251_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg365_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg330_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg127_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add3_0_impl_0_out);

   Delay1No60_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_0_impl_0_out,
                 Y => Delay1No60_out);

SharedReg301_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg301_out;
SharedReg18_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg18_out;
SharedReg24_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg24_out;
SharedReg328_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg328_out;
SharedReg480_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg480_out;
SharedReg850_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg850_out;
SharedReg334_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg334_out;
SharedReg297_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg297_out;
SharedReg363_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg363_out;
SharedReg250_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg250_out;
SharedReg849_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg849_out;
SharedReg624_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg624_out;
   MUX_Add3_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg301_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg18_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg849_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg624_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg24_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg328_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg480_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg850_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg334_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg297_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg363_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg250_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add3_0_impl_1_out);

   Delay1No61_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_0_impl_1_out,
                 Y => Delay1No61_out);

Delay1No62_out_to_Add3_1_impl_parent_implementedSystem_port_0_cast <= Delay1No62_out;
Delay1No63_out_to_Add3_1_impl_parent_implementedSystem_port_1_cast <= Delay1No63_out;
   Add3_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add3_1_impl_out,
                 X => Delay1No62_out_to_Add3_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No63_out_to_Add3_1_impl_parent_implementedSystem_port_1_cast);

SharedReg235_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg235_out;
SharedReg484_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg484_out;
SharedReg375_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg375_out;
SharedReg2_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg2_out;
SharedReg8_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg8_out;
SharedReg419_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg419_out;
SharedReg552_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg552_out;
SharedReg254_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg254_out;
SharedReg1044_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1044_out;
SharedReg40_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg40_out;
SharedReg373_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg373_out;
SharedReg130_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg130_out;
   MUX_Add3_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg235_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg484_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg373_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg130_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg375_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg2_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg8_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg419_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg552_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg254_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1044_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg40_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add3_1_impl_0_out);

   Delay1No62_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_1_impl_0_out,
                 Y => Delay1No62_out);

SharedReg372_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg372_out;
SharedReg627_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg627_out;
SharedReg259_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg259_out;
SharedReg18_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg18_out;
SharedReg24_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg24_out;
SharedReg484_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg484_out;
SharedReg606_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg606_out;
SharedReg131_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg131_out;
SharedReg574_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg574_out;
SharedReg164_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg164_out;
SharedReg164_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg164_out;
SharedReg336_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg336_out;
   MUX_Add3_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg372_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg627_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg164_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg336_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg259_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg18_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg24_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg484_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg606_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg131_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg574_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg164_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add3_1_impl_1_out);

   Delay1No63_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_1_impl_1_out,
                 Y => Delay1No63_out);

Delay1No64_out_to_Add3_2_impl_parent_implementedSystem_port_0_cast <= Delay1No64_out;
Delay1No65_out_to_Add3_2_impl_parent_implementedSystem_port_1_cast <= Delay1No65_out;
   Add3_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add3_2_impl_out,
                 X => Delay1No64_out_to_Add3_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No65_out_to_Add3_2_impl_parent_implementedSystem_port_1_cast);

SharedReg343_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg343_out;
SharedReg105_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg105_out;
SharedReg577_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg577_out;
SharedReg509_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg509_out;
SharedReg682_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg682_out;
SharedReg2_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg2_out;
SharedReg8_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg8_out;
SharedReg421_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg421_out;
SharedReg554_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg554_out;
SharedReg302_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg302_out;
SharedReg1049_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1049_out;
SharedReg76_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg76_out;
   MUX_Add3_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg343_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg105_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1049_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg76_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg577_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg509_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg682_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg2_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg8_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg421_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg554_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg302_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add3_2_impl_0_out);

   Delay1No64_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_2_impl_0_out,
                 Y => Delay1No64_out);

SharedReg170_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg170_out;
SharedReg240_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg240_out;
SharedReg576_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg576_out;
SharedReg535_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg535_out;
SharedReg789_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg789_out;
SharedReg18_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg18_out;
SharedReg24_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg24_out;
SharedReg487_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg487_out;
SharedReg609_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg609_out;
SharedReg240_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg240_out;
SharedReg449_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg449_out;
SharedReg170_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg170_out;
   MUX_Add3_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg170_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg240_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg449_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg170_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg576_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg535_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg789_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg18_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg24_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg487_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg609_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg240_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add3_2_impl_1_out);

   Delay1No65_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_2_impl_1_out,
                 Y => Delay1No65_out);

Delay1No66_out_to_Add3_3_impl_parent_implementedSystem_port_0_cast <= Delay1No66_out;
Delay1No67_out_to_Add3_3_impl_parent_implementedSystem_port_1_cast <= Delay1No67_out;
   Add3_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add3_3_impl_out,
                 X => Delay1No66_out_to_Add3_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No67_out_to_Add3_3_impl_parent_implementedSystem_port_1_cast);

SharedReg582_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg582_out;
SharedReg351_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg351_out;
SharedReg110_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg110_out;
SharedReg581_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg581_out;
SharedReg490_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg490_out;
SharedReg195_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg195_out;
SharedReg2_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg2_out;
SharedReg9_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg9_out;
SharedReg423_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg423_out;
SharedReg730_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg730_out;
SharedReg456_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg456_out;
SharedReg352_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg352_out;
   MUX_Add3_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg582_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg351_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg456_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg352_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg110_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg581_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg490_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg195_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg2_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg9_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg423_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg730_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add3_3_impl_0_out);

   Delay1No66_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_3_impl_0_out,
                 Y => Delay1No66_out);

SharedReg580_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg580_out;
SharedReg175_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg175_out;
SharedReg351_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg351_out;
SharedReg580_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg580_out;
SharedReg633_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg633_out;
SharedReg248_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg248_out;
SharedReg18_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg18_out;
SharedReg25_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg25_out;
SharedReg490_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg490_out;
SharedReg809_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg809_out;
SharedReg991_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg991_out;
SharedReg354_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg354_out;
   MUX_Add3_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg580_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg175_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg991_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg354_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg351_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg580_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg633_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg248_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg18_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg25_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg490_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg809_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add3_3_impl_1_out);

   Delay1No67_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_3_impl_1_out,
                 Y => Delay1No67_out);

Delay1No68_out_to_Add3_4_impl_parent_implementedSystem_port_0_cast <= Delay1No68_out;
Delay1No69_out_to_Add3_4_impl_parent_implementedSystem_port_1_cast <= Delay1No69_out;
   Add3_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add3_4_impl_out,
                 X => Delay1No68_out_to_Add3_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No69_out_to_Add3_4_impl_parent_implementedSystem_port_1_cast);

SharedReg709_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg709_out;
SharedReg797_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg797_out;
SharedReg84_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg84_out;
SharedReg282_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg282_out;
SharedReg81_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg81_out;
SharedReg459_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg459_out;
SharedReg517_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg517_out;
SharedReg283_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg283_out;
SharedReg2_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg2_out;
SharedReg9_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg9_out;
Delay6No4_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_11_cast <= Delay6No4_out;
SharedReg734_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg734_out;
   MUX_Add3_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg709_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg797_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay6No4_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg734_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg84_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg282_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg81_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg459_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg517_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg283_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg2_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg9_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add3_4_impl_0_out);

   Delay1No68_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_4_impl_0_out,
                 Y => Delay1No68_out);

SharedReg994_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg994_out;
SharedReg463_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg463_out;
SharedReg278_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg278_out;
SharedReg308_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg308_out;
SharedReg146_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg146_out;
SharedReg458_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg458_out;
SharedReg541_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg541_out;
SharedReg277_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg277_out;
SharedReg18_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg18_out;
SharedReg25_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg25_out;
SharedReg519_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg519_out;
SharedReg812_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg812_out;
   MUX_Add3_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg994_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg463_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg519_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg812_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg278_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg308_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg146_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg458_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg541_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg277_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg18_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg25_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add3_4_impl_1_out);

   Delay1No69_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_4_impl_1_out,
                 Y => Delay1No69_out);

Delay1No70_out_to_Add3_5_impl_parent_implementedSystem_port_0_cast <= Delay1No70_out;
Delay1No71_out_to_Add3_5_impl_parent_implementedSystem_port_1_cast <= Delay1No71_out;
   Add3_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add3_5_impl_out,
                 X => Delay1No70_out_to_Add3_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No71_out_to_Add3_5_impl_parent_implementedSystem_port_1_cast);

SharedReg427_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg427_out;
SharedReg426_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg426_out;
SharedReg712_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg712_out;
SharedReg1030_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1030_out;
SharedReg773_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg773_out;
SharedReg715_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg715_out;
SharedReg464_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg464_out;
SharedReg119_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg119_out;
SharedReg410_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg410_out;
SharedReg592_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg592_out;
SharedReg2_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg2_out;
SharedReg8_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg8_out;
   MUX_Add3_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg427_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg426_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg2_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg8_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg712_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1030_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg773_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg715_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg464_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg119_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg410_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg592_out_to_MUX_Add3_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add3_5_impl_0_out);

   Delay1No70_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_5_impl_0_out,
                 Y => Delay1No70_out);

SharedReg496_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg496_out;
SharedReg495_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg495_out;
SharedReg869_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg869_out;
SharedReg472_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg472_out;
SharedReg764_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg764_out;
SharedReg868_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg868_out;
SharedReg590_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg590_out;
SharedReg286_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg286_out;
SharedReg427_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg427_out;
SharedReg717_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg717_out;
SharedReg18_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg18_out;
SharedReg24_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg24_out;
   MUX_Add3_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg496_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg495_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg18_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg24_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg869_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg472_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg764_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg868_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg590_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg286_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg427_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg717_out_to_MUX_Add3_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add3_5_impl_1_out);

   Delay1No71_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_5_impl_1_out,
                 Y => Delay1No71_out);

Delay1No72_out_to_Add3_6_impl_parent_implementedSystem_port_0_cast <= Delay1No72_out;
Delay1No73_out_to_Add3_6_impl_parent_implementedSystem_port_1_cast <= Delay1No73_out;
   Add3_6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add3_6_impl_out,
                 X => Delay1No72_out_to_Add3_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No73_out_to_Add3_6_impl_parent_implementedSystem_port_1_cast);

SharedReg9_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg9_out;
SharedReg323_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg323_out;
SharedReg562_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg562_out;
SharedReg473_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg473_out;
SharedReg220_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg220_out;
SharedReg384_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg384_out;
SharedReg599_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg599_out;
SharedReg123_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg123_out;
SharedReg92_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg92_out;
SharedReg499_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg499_out;
SharedReg359_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg359_out;
SharedReg2_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg2_out;
   MUX_Add3_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg9_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg323_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg359_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg2_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg562_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg473_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg220_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg384_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg599_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg123_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg92_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg499_out_to_MUX_Add3_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add3_6_impl_0_out);

   Delay1No72_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_6_impl_0_out,
                 Y => Delay1No72_out);

SharedReg25_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg25_out;
SharedReg383_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg383_out;
SharedReg621_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg621_out;
SharedReg872_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg872_out;
SharedReg362_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg362_out;
SharedReg218_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg218_out;
SharedReg1066_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1066_out;
SharedReg219_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg219_out;
SharedReg320_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg320_out;
SharedReg642_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg642_out;
SharedReg325_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg325_out;
SharedReg18_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg18_out;
   MUX_Add3_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg25_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg383_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg325_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg18_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg621_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg872_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg362_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg218_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1066_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg219_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg320_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg642_out_to_MUX_Add3_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add3_6_impl_1_out);

   Delay1No73_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_6_impl_1_out,
                 Y => Delay1No73_out);

Delay1No74_out_to_Add12_0_impl_parent_implementedSystem_port_0_cast <= Delay1No74_out;
Delay1No75_out_to_Add12_0_impl_parent_implementedSystem_port_1_cast <= Delay1No75_out;
   Add12_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add12_0_impl_out,
                 X => Delay1No74_out_to_Add12_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No75_out_to_Add12_0_impl_parent_implementedSystem_port_1_cast);

SharedReg852_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg852_out;
SharedReg3_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg3_out;
SharedReg9_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg9_out;
SharedReg417_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg417_out;
SharedReg550_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg550_out;
SharedReg249_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg249_out;
SharedReg1039_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1039_out;
SharedReg35_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg35_out;
SharedReg327_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg327_out;
SharedReg202_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg202_out;
SharedReg250_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg250_out;
SharedReg551_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg551_out;
   MUX_Add12_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg852_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg3_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg250_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg551_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg9_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg417_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg550_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg249_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1039_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg35_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg327_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg202_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add12_0_impl_0_out);

   Delay1No74_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_0_impl_0_out,
                 Y => Delay1No74_out);

SharedReg671_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg671_out;
SharedReg19_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg19_out;
SharedReg25_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg25_out;
SharedReg481_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg481_out;
SharedReg603_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg603_out;
SharedReg128_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg128_out;
SharedReg670_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg670_out;
SharedReg363_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg363_out;
SharedReg158_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg158_out;
SharedReg327_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg327_out;
SharedReg363_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg363_out;
SharedReg821_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg821_out;
   MUX_Add12_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg671_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg19_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg363_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg821_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg25_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg481_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg603_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg128_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg670_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg363_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg158_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg327_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add12_0_impl_1_out);

   Delay1No75_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_0_impl_1_out,
                 Y => Delay1No75_out);

Delay1No76_out_to_Add12_1_impl_parent_implementedSystem_port_0_cast <= Delay1No76_out;
Delay1No77_out_to_Add12_1_impl_parent_implementedSystem_port_1_cast <= Delay1No77_out;
   Add12_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add12_1_impl_out,
                 X => Delay1No76_out_to_Add12_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No77_out_to_Add12_1_impl_parent_implementedSystem_port_1_cast);

SharedReg373_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg373_out;
SharedReg553_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg553_out;
SharedReg857_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg857_out;
SharedReg3_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg3_out;
SharedReg9_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg9_out;
Delay6No1_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_6_cast <= Delay6No1_out;
SharedReg722_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg722_out;
SharedReg573_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg573_out;
SharedReg337_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg337_out;
SharedReg572_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg572_out;
SharedReg675_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg675_out;
SharedReg854_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg854_out;
   MUX_Add12_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg373_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg553_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg675_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg854_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg857_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg3_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg9_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay6No1_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg722_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg573_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg337_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg572_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add12_1_impl_0_out);

   Delay1No76_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_1_impl_0_out,
                 Y => Delay1No76_out);

SharedReg340_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg340_out;
SharedReg825_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg825_out;
SharedReg575_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg575_out;
SharedReg19_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg19_out;
SharedReg25_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg25_out;
SharedReg507_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg507_out;
SharedReg803_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg803_out;
SharedReg985_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg985_out;
SharedReg379_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg379_out;
SharedReg672_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg672_out;
SharedReg775_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg775_out;
SharedReg781_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg781_out;
   MUX_Add12_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg340_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg825_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg775_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg781_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg575_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg19_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg25_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg507_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg803_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg985_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg379_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg672_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add12_1_impl_1_out);

   Delay1No77_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_1_impl_1_out,
                 Y => Delay1No77_out);

Delay1No78_out_to_Add12_2_impl_parent_implementedSystem_port_0_cast <= Delay1No78_out;
Delay1No79_out_to_Add12_2_impl_parent_implementedSystem_port_1_cast <= Delay1No79_out;
   Add12_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add12_2_impl_out,
                 X => Delay1No78_out_to_Add12_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No79_out_to_Add12_2_impl_parent_implementedSystem_port_1_cast);

SharedReg681_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg681_out;
SharedReg134_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg134_out;
SharedReg240_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg240_out;
SharedReg487_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg487_out;
SharedReg173_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg173_out;
SharedReg3_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg3_out;
SharedReg9_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg9_out;
Delay6No2_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_8_cast <= Delay6No2_out;
SharedReg726_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg726_out;
SharedReg448_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg448_out;
SharedReg344_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg344_out;
SharedReg578_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg578_out;
   MUX_Add12_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg681_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg134_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg344_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg578_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg240_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg487_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg173_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg3_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg9_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay6No2_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg726_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg448_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add12_2_impl_0_out);

   Delay1No78_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_2_impl_0_out,
                 Y => Delay1No78_out);

SharedReg783_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg783_out;
SharedReg303_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg303_out;
SharedReg342_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg342_out;
SharedReg630_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg630_out;
SharedReg265_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg265_out;
SharedReg19_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg19_out;
SharedReg25_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg25_out;
SharedReg511_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg511_out;
SharedReg806_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg806_out;
SharedReg987_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg987_out;
SharedReg348_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg348_out;
SharedReg576_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg576_out;
   MUX_Add12_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg783_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg303_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg348_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg576_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg342_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg630_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg265_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg19_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg25_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg511_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg806_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg987_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add12_2_impl_1_out);

   Delay1No79_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_2_impl_1_out,
                 Y => Delay1No79_out);

Delay1No80_out_to_Add12_3_impl_parent_implementedSystem_port_0_cast <= Delay1No80_out;
Delay1No81_out_to_Add12_3_impl_parent_implementedSystem_port_1_cast <= Delay1No81_out;
   Add12_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add12_3_impl_out,
                 X => Delay1No80_out_to_Add12_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No81_out_to_Add12_3_impl_parent_implementedSystem_port_1_cast);

SharedReg80_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg80_out;
SharedReg686_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg686_out;
SharedReg683_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg683_out;
SharedReg140_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg140_out;
SharedReg557_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg557_out;
SharedReg864_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg864_out;
SharedReg3_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg3_out;
SharedReg11_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg11_out;
Delay6No3_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_9_cast <= Delay6No3_out;
SharedReg923_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg923_out;
SharedReg422_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg422_out;
SharedReg422_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg422_out;
   MUX_Add12_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg80_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg686_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg422_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg422_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg683_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg140_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg557_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg864_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg3_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg11_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay6No3_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg923_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add12_3_impl_0_out);

   Delay1No80_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_3_impl_0_out,
                 Y => Delay1No80_out);

SharedReg175_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg175_out;
SharedReg753_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg753_out;
SharedReg881_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg881_out;
SharedReg350_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg350_out;
SharedReg833_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg833_out;
SharedReg583_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg583_out;
SharedReg19_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg19_out;
SharedReg27_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg27_out;
SharedReg515_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg515_out;
SharedReg948_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg948_out;
SharedReg489_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg489_out;
SharedReg489_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg489_out;
   MUX_Add12_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg175_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg753_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg489_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg489_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg881_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg350_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg833_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg583_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg19_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg27_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg515_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg948_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add12_3_impl_1_out);

   Delay1No81_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_3_impl_1_out,
                 Y => Delay1No81_out);

Delay1No82_out_to_Add12_4_impl_parent_implementedSystem_port_0_cast <= Delay1No82_out;
Delay1No83_out_to_Add12_4_impl_parent_implementedSystem_port_1_cast <= Delay1No83_out;
   Add12_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add12_4_impl_out,
                 X => Delay1No82_out_to_Add12_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No83_out_to_Add12_4_impl_parent_implementedSystem_port_1_cast);

SharedReg424_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg424_out;
SharedReg280_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg280_out;
SharedReg586_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg586_out;
SharedReg309_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg309_out;
SharedReg114_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg114_out;
SharedReg146_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg146_out;
SharedReg493_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg493_out;
SharedReg693_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg693_out;
SharedReg3_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg3_out;
SharedReg11_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg11_out;
SharedReg559_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg559_out;
SharedReg927_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg927_out;
   MUX_Add12_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg424_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg280_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg559_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg927_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg586_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg309_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg114_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg146_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg493_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg693_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg3_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg11_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add12_4_impl_0_out);

   Delay1No82_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_4_impl_0_out,
                 Y => Delay1No82_out);

SharedReg492_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg492_out;
SharedReg285_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg285_out;
SharedReg458_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg458_out;
SharedReg278_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg278_out;
SharedReg273_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg273_out;
SharedReg308_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg308_out;
SharedReg636_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg636_out;
SharedReg588_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg588_out;
SharedReg19_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg19_out;
SharedReg27_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg27_out;
SharedReg616_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg616_out;
SharedReg951_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg951_out;
   MUX_Add12_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg492_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg285_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg616_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg951_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg458_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg278_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg273_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg308_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg636_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg588_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg19_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg27_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add12_4_impl_1_out);

   Delay1No83_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_4_impl_1_out,
                 Y => Delay1No83_out);

Delay1No84_out_to_Add12_5_impl_parent_implementedSystem_port_0_cast <= Delay1No84_out;
Delay1No85_out_to_Add12_5_impl_parent_implementedSystem_port_1_cast <= Delay1No85_out;
   Add12_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add12_5_impl_out,
                 X => Delay1No84_out_to_Add12_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No85_out_to_Add12_5_impl_parent_implementedSystem_port_1_cast);

Delay6No5_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_1_cast <= Delay6No5_out;
SharedReg560_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg560_out;
SharedReg286_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg286_out;
SharedReg292_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg292_out;
SharedReg63_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg63_out;
SharedReg316_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg316_out;
SharedReg712_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg712_out;
SharedReg590_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg590_out;
SharedReg521_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg521_out;
SharedReg317_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg317_out;
SharedReg3_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg3_out;
SharedReg9_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg9_out;
   MUX_Add12_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay6No5_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg560_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg3_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg9_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg286_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg292_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg63_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg316_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg712_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg590_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg521_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg317_out_to_MUX_Add12_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add12_5_impl_0_out);

   Delay1No84_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_5_impl_0_out,
                 Y => Delay1No84_out);

SharedReg523_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg523_out;
SharedReg618_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg618_out;
SharedReg213_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg213_out;
SharedReg319_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg319_out;
SharedReg286_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg286_out;
SharedReg290_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg290_out;
SharedReg713_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg713_out;
SharedReg589_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg589_out;
SharedReg544_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg544_out;
SharedReg296_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg296_out;
SharedReg19_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg19_out;
SharedReg25_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg25_out;
   MUX_Add12_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg523_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg618_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg19_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg25_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg213_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg319_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg286_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg290_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg713_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg589_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg544_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg296_out_to_MUX_Add12_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add12_5_impl_1_out);

   Delay1No85_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_5_impl_1_out,
                 Y => Delay1No85_out);

Delay1No86_out_to_Add12_6_impl_parent_implementedSystem_port_0_cast <= Delay1No86_out;
Delay1No87_out_to_Add12_6_impl_parent_implementedSystem_port_1_cast <= Delay1No87_out;
   Add12_6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add12_6_impl_out,
                 X => Delay1No86_out_to_Add12_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No87_out_to_Add12_6_impl_parent_implementedSystem_port_1_cast);

SharedReg11_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg11_out;
SharedReg429_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg429_out;
SharedReg742_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg742_out;
SharedReg218_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg218_out;
SharedReg1068_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1068_out;
SharedReg63_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg63_out;
SharedReg385_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg385_out;
SharedReg153_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg153_out;
SharedReg700_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg700_out;
SharedReg563_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg563_out;
SharedReg873_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg873_out;
SharedReg3_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg3_out;
   MUX_Add12_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg11_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg429_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg873_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg3_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg742_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg218_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1068_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg63_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg385_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg153_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg700_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg563_out_to_MUX_Add12_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add12_6_impl_0_out);

   Delay1No86_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_6_impl_0_out,
                 Y => Delay1No86_out);

SharedReg27_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg27_out;
SharedReg499_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg499_out;
SharedReg818_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg818_out;
SharedReg154_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg154_out;
SharedReg704_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg704_out;
SharedReg355_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg355_out;
SharedReg381_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg381_out;
SharedReg356_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg356_out;
SharedReg871_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg871_out;
SharedReg845_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg845_out;
SharedReg875_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg875_out;
SharedReg19_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg19_out;
   MUX_Add12_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg27_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg499_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg875_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg19_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg818_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg154_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg704_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg355_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg381_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg356_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg871_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg845_out_to_MUX_Add12_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add12_6_impl_1_out);

   Delay1No87_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_6_impl_1_out,
                 Y => Delay1No87_out);

Delay1No88_out_to_Add5_1_impl_parent_implementedSystem_port_0_cast <= Delay1No88_out;
Delay1No89_out_to_Add5_1_impl_parent_implementedSystem_port_1_cast <= Delay1No89_out;
   Add5_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add5_1_impl_out,
                 X => Delay1No88_out_to_Add5_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No89_out_to_Add5_1_impl_parent_implementedSystem_port_1_cast);

SharedReg776_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg776_out;
SharedReg15_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg15_out;
SharedReg719_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg719_out;
SharedReg962_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg962_out;
SharedReg912_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg912_out;
SharedReg442_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg442_out;
SharedReg780_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg780_out;
SharedReg1007_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1007_out;
SharedReg339_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg339_out;
SharedReg570_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg570_out;
SharedReg103_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg103_out;
SharedReg570_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg570_out;
   MUX_Add5_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg776_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg15_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg103_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg570_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg719_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg962_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg912_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg442_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg780_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1007_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg339_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg570_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add5_1_impl_0_out);

   Delay1No88_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add5_1_impl_0_out,
                 Y => Delay1No88_out);

SharedReg438_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg438_out;
SharedReg31_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg31_out;
SharedReg801_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg801_out;
SharedReg914_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg914_out;
SharedReg940_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg940_out;
SharedReg777_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg777_out;
SharedReg777_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg777_out;
SharedReg570_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg570_out;
SharedReg236_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg236_out;
SharedReg854_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg854_out;
SharedReg130_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg130_out;
SharedReg855_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg855_out;
   MUX_Add5_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg438_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg31_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg130_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg855_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg801_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg914_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg940_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg777_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg777_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg570_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg236_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg854_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add5_1_impl_1_out);

   Delay1No89_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add5_1_impl_1_out,
                 Y => Delay1No89_out);

Delay1No90_out_to_Add5_2_impl_parent_implementedSystem_port_0_cast <= Delay1No90_out;
Delay1No91_out_to_Add5_2_impl_parent_implementedSystem_port_1_cast <= Delay1No91_out;
   Add5_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add5_2_impl_out,
                 X => Delay1No90_out_to_Add5_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No91_out_to_Add5_2_impl_parent_implementedSystem_port_1_cast);

SharedReg137_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg137_out;
SharedReg964_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg964_out;
SharedReg918_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg918_out;
SharedReg13_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg13_out;
SharedReg827_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg827_out;
SharedReg965_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg965_out;
SharedReg916_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg916_out;
SharedReg750_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg750_out;
SharedReg787_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg787_out;
SharedReg1012_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1012_out;
SharedReg305_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg305_out;
SharedReg445_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg445_out;
   MUX_Add5_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg137_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg964_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg305_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg445_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg918_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg13_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg827_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg965_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg916_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg750_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg787_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1012_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add5_2_impl_0_out);

   Delay1No90_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add5_2_impl_0_out,
                 Y => Delay1No90_out);

SharedReg134_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg134_out;
SharedReg942_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg942_out;
Delay4No260_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_3_cast <= Delay4No260_out;
SharedReg29_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg29_out;
SharedReg628_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg628_out;
SharedReg918_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg918_out;
SharedReg943_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg943_out;
SharedReg785_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg785_out;
SharedReg747_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg747_out;
SharedReg576_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg576_out;
SharedReg262_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg262_out;
SharedReg678_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg678_out;
   MUX_Add5_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg134_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg942_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg262_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg678_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => Delay4No260_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg29_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg628_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg918_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg943_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg785_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg747_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg576_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add5_2_impl_1_out);

   Delay1No91_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add5_2_impl_1_out,
                 Y => Delay1No91_out);

Delay1No92_out_to_Add5_3_impl_parent_implementedSystem_port_0_cast <= Delay1No92_out;
Delay1No93_out_to_Add5_3_impl_parent_implementedSystem_port_1_cast <= Delay1No93_out;
   Add5_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add5_3_impl_out,
                 X => Delay1No92_out_to_Add5_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No93_out_to_Add5_3_impl_parent_implementedSystem_port_1_cast);

SharedReg451_out_to_MUX_Add5_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg451_out;
SharedReg986_out_to_MUX_Add5_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg986_out;
SharedReg632_out_to_MUX_Add5_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg632_out;
SharedReg919_out_to_MUX_Add5_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg919_out;
Delay4No219_out_to_MUX_Add5_3_impl_0_parent_implementedSystem_port_5_cast <= Delay4No219_out;
SharedReg13_out_to_MUX_Add5_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg13_out;
SharedReg831_out_to_MUX_Add5_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg831_out;
SharedReg968_out_to_MUX_Add5_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg968_out;
SharedReg920_out_to_MUX_Add5_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg920_out;
SharedReg880_out_to_MUX_Add5_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg880_out;
SharedReg1017_out_to_MUX_Add5_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1017_out;
SharedReg269_out_to_MUX_Add5_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg269_out;
   MUX_Add5_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg451_out_to_MUX_Add5_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg986_out_to_MUX_Add5_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1017_out_to_MUX_Add5_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg269_out_to_MUX_Add5_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg632_out_to_MUX_Add5_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg919_out_to_MUX_Add5_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay4No219_out_to_MUX_Add5_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg13_out_to_MUX_Add5_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg831_out_to_MUX_Add5_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg968_out_to_MUX_Add5_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg920_out_to_MUX_Add5_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg880_out_to_MUX_Add5_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add5_3_impl_0_out);

   Delay1No92_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add5_3_impl_0_out,
                 Y => Delay1No92_out);

SharedReg683_out_to_MUX_Add5_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg683_out;
SharedReg989_out_to_MUX_Add5_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg989_out;
SharedReg403_out_to_MUX_Add5_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg403_out;
SharedReg892_out_to_MUX_Add5_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg892_out;
Delay4No226_out_to_MUX_Add5_3_impl_1_parent_implementedSystem_port_5_cast <= Delay4No226_out;
SharedReg29_out_to_MUX_Add5_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg29_out;
SharedReg631_out_to_MUX_Add5_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg631_out;
SharedReg922_out_to_MUX_Add5_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg922_out;
SharedReg946_out_to_MUX_Add5_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg946_out;
SharedReg755_out_to_MUX_Add5_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg755_out;
SharedReg580_out_to_MUX_Add5_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg580_out;
SharedReg246_out_to_MUX_Add5_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg246_out;
   MUX_Add5_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg683_out_to_MUX_Add5_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg989_out_to_MUX_Add5_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg580_out_to_MUX_Add5_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg246_out_to_MUX_Add5_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg403_out_to_MUX_Add5_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg892_out_to_MUX_Add5_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay4No226_out_to_MUX_Add5_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg29_out_to_MUX_Add5_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg631_out_to_MUX_Add5_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg922_out_to_MUX_Add5_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg946_out_to_MUX_Add5_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg755_out_to_MUX_Add5_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add5_3_impl_1_out);

   Delay1No93_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add5_3_impl_1_out,
                 Y => Delay1No93_out);

Delay1No94_out_to_Add5_4_impl_parent_implementedSystem_port_0_cast <= Delay1No94_out;
Delay1No95_out_to_Add5_4_impl_parent_implementedSystem_port_1_cast <= Delay1No95_out;
   Add5_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add5_4_impl_out,
                 X => Delay1No94_out_to_Add5_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No95_out_to_Add5_4_impl_parent_implementedSystem_port_1_cast);

SharedReg53_out_to_MUX_Add5_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg53_out;
SharedReg275_out_to_MUX_Add5_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg275_out;
SharedReg705_out_to_MUX_Add5_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg705_out;
SharedReg635_out_to_MUX_Add5_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg635_out;
SharedReg970_out_to_MUX_Add5_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg970_out;
SharedReg926_out_to_MUX_Add5_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg926_out;
SharedReg13_out_to_MUX_Add5_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg13_out;
SharedReg731_out_to_MUX_Add5_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg731_out;
SharedReg971_out_to_MUX_Add5_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg971_out;
SharedReg12_out_to_MUX_Add5_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg12_out;
SharedReg85_out_to_MUX_Add5_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg85_out;
SharedReg462_out_to_MUX_Add5_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg462_out;
   MUX_Add5_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg53_out_to_MUX_Add5_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg275_out_to_MUX_Add5_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg85_out_to_MUX_Add5_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg462_out_to_MUX_Add5_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg705_out_to_MUX_Add5_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg635_out_to_MUX_Add5_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg970_out_to_MUX_Add5_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg926_out_to_MUX_Add5_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg13_out_to_MUX_Add5_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg731_out_to_MUX_Add5_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg971_out_to_MUX_Add5_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg12_out_to_MUX_Add5_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add5_4_impl_0_out);

   Delay1No94_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add5_4_impl_0_out,
                 Y => Delay1No94_out);

SharedReg308_out_to_MUX_Add5_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg308_out;
SharedReg274_out_to_MUX_Add5_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg274_out;
SharedReg584_out_to_MUX_Add5_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg584_out;
SharedReg406_out_to_MUX_Add5_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg406_out;
SharedReg948_out_to_MUX_Add5_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg948_out;
Delay4No262_out_to_MUX_Add5_4_impl_1_parent_implementedSystem_port_6_cast <= Delay4No262_out;
SharedReg29_out_to_MUX_Add5_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg29_out;
SharedReg810_out_to_MUX_Add5_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg810_out;
SharedReg926_out_to_MUX_Add5_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg926_out;
SharedReg28_out_to_MUX_Add5_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg28_out;
SharedReg310_out_to_MUX_Add5_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg310_out;
SharedReg460_out_to_MUX_Add5_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg460_out;
   MUX_Add5_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg308_out_to_MUX_Add5_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg274_out_to_MUX_Add5_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg310_out_to_MUX_Add5_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg460_out_to_MUX_Add5_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg584_out_to_MUX_Add5_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg406_out_to_MUX_Add5_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg948_out_to_MUX_Add5_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay4No262_out_to_MUX_Add5_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg29_out_to_MUX_Add5_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg810_out_to_MUX_Add5_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg926_out_to_MUX_Add5_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg28_out_to_MUX_Add5_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add5_4_impl_1_out);

   Delay1No95_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add5_4_impl_1_out,
                 Y => Delay1No95_out);

Delay1No96_out_to_Add14_5_impl_parent_implementedSystem_port_0_cast <= Delay1No96_out;
Delay1No97_out_to_Add14_5_impl_parent_implementedSystem_port_1_cast <= Delay1No97_out;
   Add14_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add14_5_impl_out,
                 X => Delay1No96_out_to_Add14_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No97_out_to_Add14_5_impl_parent_implementedSystem_port_1_cast);

SharedReg561_out_to_MUX_Add14_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg561_out;
SharedReg738_out_to_MUX_Add14_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg738_out;
SharedReg469_out_to_MUX_Add14_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg469_out;
SharedReg1061_out_to_MUX_Add14_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1061_out;
SharedReg121_out_to_MUX_Add14_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg121_out;
SharedReg291_out_to_MUX_Add14_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg291_out;
SharedReg150_out_to_MUX_Add14_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg150_out;
SharedReg213_out_to_MUX_Add14_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg213_out;
SharedReg496_out_to_MUX_Add14_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg496_out;
SharedReg698_out_to_MUX_Add14_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg698_out;
SharedReg4_out_to_MUX_Add14_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg4_out;
SharedReg11_out_to_MUX_Add14_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg11_out;
   MUX_Add14_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg561_out_to_MUX_Add14_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg738_out_to_MUX_Add14_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg4_out_to_MUX_Add14_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg11_out_to_MUX_Add14_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg469_out_to_MUX_Add14_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1061_out_to_MUX_Add14_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg121_out_to_MUX_Add14_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg291_out_to_MUX_Add14_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg150_out_to_MUX_Add14_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg213_out_to_MUX_Add14_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg496_out_to_MUX_Add14_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg698_out_to_MUX_Add14_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add14_5_impl_0_out);

   Delay1No96_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add14_5_impl_0_out,
                 Y => Delay1No96_out);

SharedReg619_out_to_MUX_Add14_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg619_out;
SharedReg815_out_to_MUX_Add14_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg815_out;
SharedReg998_out_to_MUX_Add14_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg998_out;
SharedReg593_out_to_MUX_Add14_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg593_out;
SharedReg313_out_to_MUX_Add14_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg313_out;
SharedReg313_out_to_MUX_Add14_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg313_out;
SharedReg183_out_to_MUX_Add14_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg183_out;
SharedReg313_out_to_MUX_Add14_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg313_out;
SharedReg639_out_to_MUX_Add14_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg639_out;
SharedReg594_out_to_MUX_Add14_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg594_out;
SharedReg20_out_to_MUX_Add14_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg20_out;
SharedReg27_out_to_MUX_Add14_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg27_out;
   MUX_Add14_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg619_out_to_MUX_Add14_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg815_out_to_MUX_Add14_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg20_out_to_MUX_Add14_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg27_out_to_MUX_Add14_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg998_out_to_MUX_Add14_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg593_out_to_MUX_Add14_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg313_out_to_MUX_Add14_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg313_out_to_MUX_Add14_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg183_out_to_MUX_Add14_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg313_out_to_MUX_Add14_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg639_out_to_MUX_Add14_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg594_out_to_MUX_Add14_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add14_5_impl_1_out);

   Delay1No97_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add14_5_impl_1_out,
                 Y => Delay1No97_out);

Delay1No98_out_to_Add14_6_impl_parent_implementedSystem_port_0_cast <= Delay1No98_out;
Delay1No99_out_to_Add14_6_impl_parent_implementedSystem_port_1_cast <= Delay1No99_out;
   Add14_6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add14_6_impl_out,
                 X => Delay1No98_out_to_Add14_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No99_out_to_Add14_6_impl_parent_implementedSystem_port_1_cast);

SharedReg14_out_to_MUX_Add14_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg14_out;
Delay6No6_out_to_MUX_Add14_6_impl_0_parent_implementedSystem_port_2_cast <= Delay6No6_out;
SharedReg935_out_to_MUX_Add14_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg935_out;
SharedReg703_out_to_MUX_Add14_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg703_out;
SharedReg322_out_to_MUX_Add14_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg322_out;
SharedReg598_out_to_MUX_Add14_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg598_out;
SharedReg321_out_to_MUX_Add14_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg321_out;
SharedReg871_out_to_MUX_Add14_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg871_out;
SharedReg188_out_to_MUX_Add14_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg188_out;
SharedReg745_out_to_MUX_Add14_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg745_out;
SharedReg386_out_to_MUX_Add14_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg386_out;
SharedReg4_out_to_MUX_Add14_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg4_out;
   MUX_Add14_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg14_out_to_MUX_Add14_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay6No6_out_to_MUX_Add14_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg386_out_to_MUX_Add14_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg4_out_to_MUX_Add14_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg935_out_to_MUX_Add14_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg703_out_to_MUX_Add14_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg322_out_to_MUX_Add14_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg598_out_to_MUX_Add14_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg321_out_to_MUX_Add14_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg871_out_to_MUX_Add14_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg188_out_to_MUX_Add14_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg745_out_to_MUX_Add14_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add14_6_impl_0_out);

   Delay1No98_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add14_6_impl_0_out,
                 Y => Delay1No98_out);

SharedReg30_out_to_MUX_Add14_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg30_out;
SharedReg527_out_to_MUX_Add14_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg527_out;
SharedReg957_out_to_MUX_Add14_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg957_out;
SharedReg1002_out_to_MUX_Add14_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1002_out;
SharedReg388_out_to_MUX_Add14_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg388_out;
SharedReg595_out_to_MUX_Add14_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg595_out;
SharedReg389_out_to_MUX_Add14_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg389_out;
SharedReg478_out_to_MUX_Add14_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg478_out;
SharedReg381_out_to_MUX_Add14_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg381_out;
Delay4No188_out_to_MUX_Add14_6_impl_1_parent_implementedSystem_port_10_cast <= Delay4No188_out;
SharedReg394_out_to_MUX_Add14_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg394_out;
SharedReg20_out_to_MUX_Add14_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg20_out;
   MUX_Add14_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg30_out_to_MUX_Add14_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg527_out_to_MUX_Add14_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg394_out_to_MUX_Add14_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg20_out_to_MUX_Add14_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg957_out_to_MUX_Add14_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1002_out_to_MUX_Add14_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg388_out_to_MUX_Add14_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg595_out_to_MUX_Add14_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg389_out_to_MUX_Add14_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg478_out_to_MUX_Add14_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg381_out_to_MUX_Add14_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay4No188_out_to_MUX_Add14_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add14_6_impl_1_out);

   Delay1No99_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add14_6_impl_1_out,
                 Y => Delay1No99_out);

Delay1No100_out_to_Add6_4_impl_parent_implementedSystem_port_0_cast <= Delay1No100_out;
Delay1No101_out_to_Add6_4_impl_parent_implementedSystem_port_1_cast <= Delay1No101_out;
   Add6_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add6_4_impl_out,
                 X => Delay1No100_out_to_Add6_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No101_out_to_Add6_4_impl_parent_implementedSystem_port_1_cast);

SharedReg993_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg993_out;
SharedReg924_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg924_out;
SharedReg990_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg990_out;
SharedReg654_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg654_out;
SharedReg923_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg923_out;
Delay4No220_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_6_cast <= Delay4No220_out;
SharedReg10_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg10_out;
SharedReg835_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg835_out;
Delay6No45_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_9_cast <= Delay6No45_out;
SharedReg924_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg924_out;
SharedReg761_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg761_out;
SharedReg794_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg794_out;
   MUX_Add6_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg993_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg924_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg761_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg794_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg990_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg654_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg923_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay4No220_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg10_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg835_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay6No45_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg924_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add6_4_impl_0_out);

   Delay1No100_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add6_4_impl_0_out,
                 Y => Delay1No100_out);

SharedReg458_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg458_out;
SharedReg949_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg949_out;
SharedReg992_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg992_out;
SharedReg730_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg730_out;
SharedReg896_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg896_out;
Delay4No227_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_6_cast <= Delay4No227_out;
SharedReg26_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg26_out;
SharedReg634_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg634_out;
SharedReg925_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg925_out;
SharedReg949_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg949_out;
SharedReg707_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg707_out;
SharedReg707_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg707_out;
   MUX_Add6_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg458_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg949_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg707_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg707_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg992_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg730_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg896_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay4No227_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg26_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg634_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg925_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg949_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add6_4_impl_1_out);

   Delay1No101_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add6_4_impl_1_out,
                 Y => Delay1No101_out);

Delay1No102_out_to_Add15_3_impl_parent_implementedSystem_port_0_cast <= Delay1No102_out;
Delay1No103_out_to_Add15_3_impl_parent_implementedSystem_port_1_cast <= Delay1No103_out;
   Add15_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add15_3_impl_out,
                 X => Delay1No102_out_to_Add15_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No103_out_to_Add15_3_impl_parent_implementedSystem_port_1_cast);

SharedReg793_out_to_MUX_Add15_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg793_out;
SharedReg112_out_to_MUX_Add15_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg112_out;
SharedReg451_out_to_MUX_Add15_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg451_out;
SharedReg967_out_to_MUX_Add15_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg967_out;
SharedReg922_out_to_MUX_Add15_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg922_out;
SharedReg15_out_to_MUX_Add15_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg15_out;
SharedReg727_out_to_MUX_Add15_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg727_out;
SharedReg12_out_to_MUX_Add15_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg12_out;
SharedReg456_out_to_MUX_Add15_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg456_out;
SharedReg688_out_to_MUX_Add15_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg688_out;
SharedReg192_out_to_MUX_Add15_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg192_out;
SharedReg1019_out_to_MUX_Add15_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1019_out;
   MUX_Add15_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg793_out_to_MUX_Add15_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg112_out_to_MUX_Add15_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg192_out_to_MUX_Add15_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1019_out_to_MUX_Add15_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg451_out_to_MUX_Add15_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg967_out_to_MUX_Add15_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg922_out_to_MUX_Add15_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg15_out_to_MUX_Add15_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg727_out_to_MUX_Add15_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg12_out_to_MUX_Add15_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg456_out_to_MUX_Add15_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg688_out_to_MUX_Add15_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add15_3_impl_0_out);

   Delay1No102_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add15_3_impl_0_out,
                 Y => Delay1No102_out);

SharedReg753_out_to_MUX_Add15_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg753_out;
SharedReg139_out_to_MUX_Add15_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg139_out;
SharedReg862_out_to_MUX_Add15_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg862_out;
SharedReg945_out_to_MUX_Add15_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg945_out;
Delay4No261_out_to_MUX_Add15_3_impl_1_parent_implementedSystem_port_5_cast <= Delay4No261_out;
SharedReg31_out_to_MUX_Add15_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg31_out;
SharedReg807_out_to_MUX_Add15_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg807_out;
SharedReg28_out_to_MUX_Add15_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg28_out;
SharedReg755_out_to_MUX_Add15_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg755_out;
SharedReg453_out_to_MUX_Add15_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg453_out;
SharedReg350_out_to_MUX_Add15_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg350_out;
SharedReg757_out_to_MUX_Add15_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg757_out;
   MUX_Add15_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg753_out_to_MUX_Add15_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg139_out_to_MUX_Add15_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg350_out_to_MUX_Add15_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg757_out_to_MUX_Add15_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg862_out_to_MUX_Add15_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg945_out_to_MUX_Add15_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay4No261_out_to_MUX_Add15_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg31_out_to_MUX_Add15_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg807_out_to_MUX_Add15_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg28_out_to_MUX_Add15_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg755_out_to_MUX_Add15_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg453_out_to_MUX_Add15_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add15_3_impl_1_out);

   Delay1No103_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add15_3_impl_1_out,
                 Y => Delay1No103_out);

Delay1No104_out_to_Add8_0_impl_parent_implementedSystem_port_0_cast <= Delay1No104_out;
Delay1No105_out_to_Add8_0_impl_parent_implementedSystem_port_1_cast <= Delay1No105_out;
   Add8_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add8_0_impl_out,
                 X => Delay1No104_out_to_Add8_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No105_out_to_Add8_0_impl_parent_implementedSystem_port_1_cast);

SharedReg366_out_to_MUX_Add8_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg366_out;
SharedReg4_out_to_MUX_Add8_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg4_out;
SharedReg11_out_to_MUX_Add8_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg11_out;
Delay6No_out_to_MUX_Add8_0_impl_0_parent_implementedSystem_port_4_cast <= Delay6No_out;
SharedReg718_out_to_MUX_Add8_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg718_out;
SharedReg669_out_to_MUX_Add8_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg669_out;
SharedReg298_out_to_MUX_Add8_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg298_out;
SharedReg566_out_to_MUX_Add8_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg566_out;
SharedReg668_out_to_MUX_Add8_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg668_out;
SharedReg981_out_to_MUX_Add8_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg981_out;
SharedReg364_out_to_MUX_Add8_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg364_out;
SharedReg721_out_to_MUX_Add8_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg721_out;
   MUX_Add8_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg366_out_to_MUX_Add8_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg4_out_to_MUX_Add8_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg364_out_to_MUX_Add8_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg721_out_to_MUX_Add8_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg11_out_to_MUX_Add8_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay6No_out_to_MUX_Add8_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg718_out_to_MUX_Add8_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg669_out_to_MUX_Add8_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg298_out_to_MUX_Add8_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg566_out_to_MUX_Add8_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg668_out_to_MUX_Add8_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg981_out_to_MUX_Add8_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add8_0_impl_0_out);

   Delay1No104_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add8_0_impl_0_out,
                 Y => Delay1No104_out);

SharedReg371_out_to_MUX_Add8_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg371_out;
SharedReg20_out_to_MUX_Add8_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg20_out;
SharedReg27_out_to_MUX_Add8_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg27_out;
SharedReg503_out_to_MUX_Add8_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg503_out;
SharedReg800_out_to_MUX_Add8_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg800_out;
SharedReg982_out_to_MUX_Add8_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg982_out;
SharedReg370_out_to_MUX_Add8_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg370_out;
SharedReg666_out_to_MUX_Add8_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg666_out;
SharedReg430_out_to_MUX_Add8_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg430_out;
SharedReg436_out_to_MUX_Add8_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg436_out;
SharedReg333_out_to_MUX_Add8_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg333_out;
Delay4No182_out_to_MUX_Add8_0_impl_1_parent_implementedSystem_port_12_cast <= Delay4No182_out;
   MUX_Add8_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg371_out_to_MUX_Add8_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg20_out_to_MUX_Add8_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg333_out_to_MUX_Add8_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay4No182_out_to_MUX_Add8_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg27_out_to_MUX_Add8_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg503_out_to_MUX_Add8_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg800_out_to_MUX_Add8_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg982_out_to_MUX_Add8_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg370_out_to_MUX_Add8_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg666_out_to_MUX_Add8_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg430_out_to_MUX_Add8_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg436_out_to_MUX_Add8_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add8_0_impl_1_out);

   Delay1No105_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add8_0_impl_1_out,
                 Y => Delay1No105_out);

Delay1No106_out_to_Add8_4_impl_parent_implementedSystem_port_0_cast <= Delay1No106_out;
Delay1No107_out_to_Add8_4_impl_parent_implementedSystem_port_1_cast <= Delay1No107_out;
   Add8_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add8_4_impl_out,
                 X => Delay1No106_out_to_Add8_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No107_out_to_Add8_4_impl_parent_implementedSystem_port_1_cast);

SharedReg558_out_to_MUX_Add8_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg558_out;
SharedReg424_out_to_MUX_Add8_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg424_out;
SharedReg116_out_to_MUX_Add8_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg116_out;
SharedReg692_out_to_MUX_Add8_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg692_out;
SharedReg584_out_to_MUX_Add8_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg584_out;
SharedReg309_out_to_MUX_Add8_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg309_out;
SharedReg559_out_to_MUX_Add8_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg559_out;
SharedReg56_out_to_MUX_Add8_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg56_out;
SharedReg4_out_to_MUX_Add8_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg4_out;
SharedReg14_out_to_MUX_Add8_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg14_out;
SharedReg735_out_to_MUX_Add8_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg735_out;
SharedReg559_out_to_MUX_Add8_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg559_out;
   MUX_Add8_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg558_out_to_MUX_Add8_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg424_out_to_MUX_Add8_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg735_out_to_MUX_Add8_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg559_out_to_MUX_Add8_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg116_out_to_MUX_Add8_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg692_out_to_MUX_Add8_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg584_out_to_MUX_Add8_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg309_out_to_MUX_Add8_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg559_out_to_MUX_Add8_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg56_out_to_MUX_Add8_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg4_out_to_MUX_Add8_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg14_out_to_MUX_Add8_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add8_4_impl_0_out);

   Delay1No106_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add8_4_impl_0_out,
                 Y => Delay1No106_out);

SharedReg615_out_to_MUX_Add8_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg615_out;
SharedReg492_out_to_MUX_Add8_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg492_out;
SharedReg52_out_to_MUX_Add8_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg52_out;
SharedReg790_out_to_MUX_Add8_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg790_out;
SharedReg762_out_to_MUX_Add8_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg762_out;
SharedReg311_out_to_MUX_Add8_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg311_out;
SharedReg837_out_to_MUX_Add8_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg837_out;
SharedReg59_out_to_MUX_Add8_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg59_out;
SharedReg20_out_to_MUX_Add8_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg20_out;
SharedReg30_out_to_MUX_Add8_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg30_out;
SharedReg813_out_to_MUX_Add8_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg813_out;
SharedReg616_out_to_MUX_Add8_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg616_out;
   MUX_Add8_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg615_out_to_MUX_Add8_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg492_out_to_MUX_Add8_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg813_out_to_MUX_Add8_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg616_out_to_MUX_Add8_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg52_out_to_MUX_Add8_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg790_out_to_MUX_Add8_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg762_out_to_MUX_Add8_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg311_out_to_MUX_Add8_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg837_out_to_MUX_Add8_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg59_out_to_MUX_Add8_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg20_out_to_MUX_Add8_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg30_out_to_MUX_Add8_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add8_4_impl_1_out);

   Delay1No107_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add8_4_impl_1_out,
                 Y => Delay1No107_out);

Delay1No108_out_to_Add8_5_impl_parent_implementedSystem_port_0_cast <= Delay1No108_out;
Delay1No109_out_to_Add8_5_impl_parent_implementedSystem_port_1_cast <= Delay1No109_out;
   Add8_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add8_5_impl_out,
                 X => Delay1No108_out_to_Add8_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No109_out_to_Add8_5_impl_parent_implementedSystem_port_1_cast);

SharedReg739_out_to_MUX_Add8_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg739_out;
SharedReg931_out_to_MUX_Add8_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg931_out;
SharedReg426_out_to_MUX_Add8_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg426_out;
SharedReg315_out_to_MUX_Add8_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg315_out;
SharedReg591_out_to_MUX_Add8_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg591_out;
SharedReg697_out_to_MUX_Add8_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg697_out;
SharedReg182_out_to_MUX_Add8_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg182_out;
SharedReg314_out_to_MUX_Add8_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg314_out;
SharedReg561_out_to_MUX_Add8_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg561_out;
SharedReg228_out_to_MUX_Add8_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg228_out;
SharedReg5_out_to_MUX_Add8_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg5_out;
SharedReg14_out_to_MUX_Add8_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg14_out;
   MUX_Add8_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg739_out_to_MUX_Add8_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg931_out_to_MUX_Add8_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg5_out_to_MUX_Add8_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg14_out_to_MUX_Add8_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg426_out_to_MUX_Add8_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg315_out_to_MUX_Add8_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg591_out_to_MUX_Add8_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg697_out_to_MUX_Add8_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg182_out_to_MUX_Add8_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg314_out_to_MUX_Add8_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg561_out_to_MUX_Add8_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg228_out_to_MUX_Add8_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add8_5_impl_0_out);

   Delay1No108_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add8_5_impl_0_out,
                 Y => Delay1No108_out);

SharedReg816_out_to_MUX_Add8_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg816_out;
SharedReg954_out_to_MUX_Add8_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg954_out;
SharedReg495_out_to_MUX_Add8_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg495_out;
SharedReg232_out_to_MUX_Add8_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg232_out;
SharedReg464_out_to_MUX_Add8_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg464_out;
SharedReg795_out_to_MUX_Add8_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg795_out;
SharedReg287_out_to_MUX_Add8_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg287_out;
SharedReg318_out_to_MUX_Add8_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg318_out;
SharedReg841_out_to_MUX_Add8_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg841_out;
SharedReg233_out_to_MUX_Add8_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg233_out;
SharedReg21_out_to_MUX_Add8_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg21_out;
SharedReg30_out_to_MUX_Add8_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg30_out;
   MUX_Add8_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg816_out_to_MUX_Add8_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg954_out_to_MUX_Add8_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg21_out_to_MUX_Add8_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg30_out_to_MUX_Add8_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg495_out_to_MUX_Add8_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg232_out_to_MUX_Add8_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg464_out_to_MUX_Add8_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg795_out_to_MUX_Add8_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg287_out_to_MUX_Add8_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg318_out_to_MUX_Add8_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg841_out_to_MUX_Add8_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg233_out_to_MUX_Add8_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add8_5_impl_1_out);

   Delay1No109_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add8_5_impl_1_out,
                 Y => Delay1No109_out);

Delay1No110_out_to_Add8_6_impl_parent_implementedSystem_port_0_cast <= Delay1No110_out;
Delay1No111_out_to_Add8_6_impl_parent_implementedSystem_port_1_cast <= Delay1No111_out;
   Add8_6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add8_6_impl_out,
                 X => Delay1No110_out_to_Add8_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No111_out_to_Add8_6_impl_parent_implementedSystem_port_1_cast);

SharedReg414_out_to_MUX_Add8_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg414_out;
SharedReg563_out_to_MUX_Add8_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg563_out;
SharedReg563_out_to_MUX_Add8_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg563_out;
SharedReg428_out_to_MUX_Add8_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg428_out;
SharedReg428_out_to_MUX_Add8_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg428_out;
SharedReg94_out_to_MUX_Add8_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg94_out;
SharedReg702_out_to_MUX_Add8_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg702_out;
SharedReg218_out_to_MUX_Add8_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg218_out;
SharedReg356_out_to_MUX_Add8_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg356_out;
Delay3No244_out_to_MUX_Add8_6_impl_0_parent_implementedSystem_port_10_cast <= Delay3No244_out;
SharedReg498_out_to_MUX_Add8_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg498_out;
SharedReg5_out_to_MUX_Add8_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg5_out;
   MUX_Add8_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg414_out_to_MUX_Add8_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg563_out_to_MUX_Add8_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg498_out_to_MUX_Add8_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg5_out_to_MUX_Add8_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg563_out_to_MUX_Add8_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg428_out_to_MUX_Add8_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg428_out_to_MUX_Add8_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg94_out_to_MUX_Add8_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg702_out_to_MUX_Add8_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg218_out_to_MUX_Add8_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg356_out_to_MUX_Add8_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay3No244_out_to_MUX_Add8_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add8_6_impl_0_out);

   Delay1No110_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add8_6_impl_0_out,
                 Y => Delay1No110_out);

SharedReg745_out_to_MUX_Add8_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg745_out;
SharedReg622_out_to_MUX_Add8_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg622_out;
SharedReg622_out_to_MUX_Add8_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg622_out;
SharedReg498_out_to_MUX_Add8_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg498_out;
SharedReg498_out_to_MUX_Add8_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg498_out;
SharedReg381_out_to_MUX_Add8_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg381_out;
SharedReg473_out_to_MUX_Add8_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg473_out;
SharedReg222_out_to_MUX_Add8_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg222_out;
SharedReg361_out_to_MUX_Add8_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg361_out;
SharedReg623_out_to_MUX_Add8_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg623_out;
SharedReg525_out_to_MUX_Add8_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg525_out;
SharedReg21_out_to_MUX_Add8_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg21_out;
   MUX_Add8_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg745_out_to_MUX_Add8_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg622_out_to_MUX_Add8_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg525_out_to_MUX_Add8_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg21_out_to_MUX_Add8_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg622_out_to_MUX_Add8_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg498_out_to_MUX_Add8_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg498_out_to_MUX_Add8_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg381_out_to_MUX_Add8_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg473_out_to_MUX_Add8_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg222_out_to_MUX_Add8_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg361_out_to_MUX_Add8_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg623_out_to_MUX_Add8_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add8_6_impl_1_out);

   Delay1No111_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add8_6_impl_1_out,
                 Y => Delay1No111_out);

Delay1No112_out_to_Add10_6_impl_parent_implementedSystem_port_0_cast <= Delay1No112_out;
Delay1No113_out_to_Add10_6_impl_parent_implementedSystem_port_1_cast <= Delay1No113_out;
   Add10_6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add10_6_impl_out,
                 X => Delay1No112_out_to_Add10_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No113_out_to_Add10_6_impl_parent_implementedSystem_port_1_cast);

SharedReg12_out_to_MUX_Add10_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg12_out;
SharedReg932_out_to_MUX_Add10_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg932_out;
SharedReg477_out_to_MUX_Add10_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg477_out;
SharedReg931_out_to_MUX_Add10_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg931_out;
SharedReg738_out_to_MUX_Add10_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg738_out;
SharedReg932_out_to_MUX_Add10_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg932_out;
SharedReg290_out_to_MUX_Add10_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg290_out;
SharedReg641_out_to_MUX_Add10_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg641_out;
SharedReg931_out_to_MUX_Add10_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg931_out;
SharedReg934_out_to_MUX_Add10_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg934_out;
SharedReg15_out_to_MUX_Add10_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg15_out;
SharedReg739_out_to_MUX_Add10_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg739_out;
   MUX_Add10_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg12_out_to_MUX_Add10_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg932_out_to_MUX_Add10_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg15_out_to_MUX_Add10_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg739_out_to_MUX_Add10_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg477_out_to_MUX_Add10_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg931_out_to_MUX_Add10_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg738_out_to_MUX_Add10_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg932_out_to_MUX_Add10_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg290_out_to_MUX_Add10_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg641_out_to_MUX_Add10_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg931_out_to_MUX_Add10_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg934_out_to_MUX_Add10_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add10_6_impl_0_out);

   Delay1No112_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add10_6_impl_0_out,
                 Y => Delay1No112_out);

SharedReg28_out_to_MUX_Add10_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg28_out;
SharedReg955_out_to_MUX_Add10_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg955_out;
SharedReg475_out_to_MUX_Add10_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg475_out;
SharedReg954_out_to_MUX_Add10_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg954_out;
SharedReg815_out_to_MUX_Add10_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg815_out;
SharedReg955_out_to_MUX_Add10_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg955_out;
SharedReg295_out_to_MUX_Add10_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg295_out;
SharedReg412_out_to_MUX_Add10_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg412_out;
SharedReg904_out_to_MUX_Add10_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg904_out;
Delay4No264_out_to_MUX_Add10_6_impl_1_parent_implementedSystem_port_10_cast <= Delay4No264_out;
SharedReg31_out_to_MUX_Add10_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg31_out;
SharedReg816_out_to_MUX_Add10_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg816_out;
   MUX_Add10_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg28_out_to_MUX_Add10_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg955_out_to_MUX_Add10_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg31_out_to_MUX_Add10_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg816_out_to_MUX_Add10_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg475_out_to_MUX_Add10_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg954_out_to_MUX_Add10_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg815_out_to_MUX_Add10_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg955_out_to_MUX_Add10_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg295_out_to_MUX_Add10_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg412_out_to_MUX_Add10_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg904_out_to_MUX_Add10_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay4No264_out_to_MUX_Add10_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add10_6_impl_1_out);

   Delay1No113_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add10_6_impl_1_out,
                 Y => Delay1No113_out);

Delay1No114_out_to_Add23_1_impl_parent_implementedSystem_port_0_cast <= Delay1No114_out;
Delay1No115_out_to_Add23_1_impl_parent_implementedSystem_port_1_cast <= Delay1No115_out;
   Add23_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add23_1_impl_out,
                 X => Delay1No114_out_to_Add23_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No115_out_to_Add23_1_impl_parent_implementedSystem_port_1_cast);

SharedReg1043_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1043_out;
SharedReg725_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg725_out;
SharedReg168_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg168_out;
SharedReg4_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg4_out;
SharedReg11_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg11_out;
SharedReg553_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg553_out;
SharedReg915_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg915_out;
SharedReg418_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg418_out;
SharedReg418_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg418_out;
SharedReg72_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg72_out;
SharedReg441_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg441_out;
SharedReg254_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg254_out;
   MUX_Add23_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1043_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg725_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg441_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg254_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg168_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg4_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg11_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg553_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg915_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg418_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg418_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg72_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add23_1_impl_0_out);

   Delay1No114_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add23_1_impl_0_out,
                 Y => Delay1No114_out);

SharedReg1046_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1046_out;
Delay4No183_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_2_cast <= Delay4No183_out;
SharedReg380_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg380_out;
SharedReg20_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg20_out;
SharedReg27_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg27_out;
SharedReg607_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg607_out;
SharedReg942_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg942_out;
SharedReg483_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg483_out;
SharedReg483_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg483_out;
SharedReg41_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg41_out;
SharedReg984_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg984_out;
SharedReg237_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg237_out;
   MUX_Add23_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1046_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay4No183_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg984_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg237_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg380_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg20_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg27_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg607_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg942_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg483_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg483_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg41_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add23_1_impl_1_out);

   Delay1No115_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add23_1_impl_1_out,
                 Y => Delay1No115_out);

Delay1No116_out_to_Add23_2_impl_parent_implementedSystem_port_0_cast <= Delay1No116_out;
Delay1No117_out_to_Add23_2_impl_parent_implementedSystem_port_1_cast <= Delay1No117_out;
   Add23_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add23_2_impl_out,
                 X => Delay1No116_out_to_Add23_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No117_out_to_Add23_2_impl_parent_implementedSystem_port_1_cast);

SharedReg447_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg447_out;
SharedReg678_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg678_out;
SharedReg343_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg343_out;
SharedReg555_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg555_out;
SharedReg860_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg860_out;
SharedReg4_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg4_out;
SharedReg11_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg11_out;
SharedReg555_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg555_out;
SharedReg919_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg919_out;
SharedReg420_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg420_out;
SharedReg420_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg420_out;
SharedReg108_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg108_out;
   MUX_Add23_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg447_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg678_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg420_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg108_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg343_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg555_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg860_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg4_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg11_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg555_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg919_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg420_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add23_2_impl_0_out);

   Delay1No116_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add23_2_impl_0_out,
                 Y => Delay1No116_out);

SharedReg858_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg858_out;
SharedReg788_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg788_out;
SharedReg306_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg306_out;
SharedReg829_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg829_out;
SharedReg450_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg450_out;
SharedReg20_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg20_out;
SharedReg27_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg27_out;
SharedReg610_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg610_out;
SharedReg945_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg945_out;
SharedReg486_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg486_out;
SharedReg486_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg486_out;
SharedReg198_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg198_out;
   MUX_Add23_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg858_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg788_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg486_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg198_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg306_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg829_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg450_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg20_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg27_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg610_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg945_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg486_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add23_2_impl_1_out);

   Delay1No117_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add23_2_impl_1_out,
                 Y => Delay1No117_out);

Delay1No118_out_to_Add23_3_impl_parent_implementedSystem_port_0_cast <= Delay1No118_out;
Delay1No119_out_to_Add23_3_impl_parent_implementedSystem_port_1_cast <= Delay1No119_out;
   Add23_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add23_3_impl_out,
                 X => Delay1No118_out_to_Add23_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No119_out_to_Add23_3_impl_parent_implementedSystem_port_1_cast);

SharedReg422_out_to_MUX_Add23_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg422_out;
SharedReg454_out_to_MUX_Add23_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg454_out;
SharedReg244_out_to_MUX_Add23_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg244_out;
SharedReg351_out_to_MUX_Add23_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg351_out;
SharedReg733_out_to_MUX_Add23_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg733_out;
SharedReg180_out_to_MUX_Add23_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg180_out;
SharedReg4_out_to_MUX_Add23_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg4_out;
SharedReg14_out_to_MUX_Add23_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg14_out;
SharedReg557_out_to_MUX_Add23_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg557_out;
SharedReg557_out_to_MUX_Add23_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg557_out;
SharedReg556_out_to_MUX_Add23_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg556_out;
SharedReg556_out_to_MUX_Add23_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg556_out;
   MUX_Add23_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg422_out_to_MUX_Add23_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg454_out_to_MUX_Add23_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg556_out_to_MUX_Add23_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg556_out_to_MUX_Add23_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg244_out_to_MUX_Add23_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg351_out_to_MUX_Add23_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg733_out_to_MUX_Add23_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg180_out_to_MUX_Add23_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg4_out_to_MUX_Add23_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg14_out_to_MUX_Add23_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg557_out_to_MUX_Add23_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg557_out_to_MUX_Add23_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add23_3_impl_0_out);

   Delay1No118_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add23_3_impl_0_out,
                 Y => Delay1No118_out);

SharedReg489_out_to_MUX_Add23_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg489_out;
SharedReg990_out_to_MUX_Add23_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg990_out;
SharedReg143_out_to_MUX_Add23_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg143_out;
SharedReg270_out_to_MUX_Add23_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg270_out;
Delay4No185_out_to_MUX_Add23_3_impl_1_parent_implementedSystem_port_5_cast <= Delay4No185_out;
SharedReg197_out_to_MUX_Add23_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg197_out;
SharedReg20_out_to_MUX_Add23_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg20_out;
SharedReg30_out_to_MUX_Add23_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg30_out;
SharedReg613_out_to_MUX_Add23_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg613_out;
SharedReg613_out_to_MUX_Add23_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg613_out;
SharedReg612_out_to_MUX_Add23_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg612_out;
SharedReg612_out_to_MUX_Add23_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg612_out;
   MUX_Add23_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg489_out_to_MUX_Add23_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg990_out_to_MUX_Add23_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg612_out_to_MUX_Add23_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg612_out_to_MUX_Add23_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg143_out_to_MUX_Add23_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg270_out_to_MUX_Add23_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay4No185_out_to_MUX_Add23_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg197_out_to_MUX_Add23_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg20_out_to_MUX_Add23_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg30_out_to_MUX_Add23_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg613_out_to_MUX_Add23_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg613_out_to_MUX_Add23_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add23_3_impl_1_out);

   Delay1No119_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add23_3_impl_1_out,
                 Y => Delay1No119_out);

Delay1No120_out_to_Add113_0_impl_parent_implementedSystem_port_0_cast <= Delay1No120_out;
Delay1No121_out_to_Add113_0_impl_parent_implementedSystem_port_1_cast <= Delay1No121_out;
   Add113_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add113_0_impl_out,
                 X => Delay1No120_out_to_Add113_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No121_out_to_Add113_0_impl_parent_implementedSystem_port_1_cast);

SharedReg480_out_to_MUX_Add113_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg480_out;
SharedReg5_out_to_MUX_Add113_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg5_out;
SharedReg14_out_to_MUX_Add113_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg14_out;
SharedReg551_out_to_MUX_Add113_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg551_out;
SharedReg911_out_to_MUX_Add113_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg911_out;
SharedReg416_out_to_MUX_Add113_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg416_out;
SharedReg416_out_to_MUX_Add113_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg416_out;
SharedReg68_out_to_MUX_Add113_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg68_out;
SharedReg433_out_to_MUX_Add113_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg433_out;
SharedReg297_out_to_MUX_Add113_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg297_out;
SharedReg1071_out_to_MUX_Add113_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1071_out;
Delay3No238_out_to_MUX_Add113_0_impl_0_parent_implementedSystem_port_12_cast <= Delay3No238_out;
   MUX_Add113_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg480_out_to_MUX_Add113_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg5_out_to_MUX_Add113_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1071_out_to_MUX_Add113_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay3No238_out_to_MUX_Add113_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg14_out_to_MUX_Add113_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg551_out_to_MUX_Add113_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg911_out_to_MUX_Add113_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg416_out_to_MUX_Add113_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg416_out_to_MUX_Add113_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg68_out_to_MUX_Add113_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg433_out_to_MUX_Add113_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg297_out_to_MUX_Add113_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add113_0_impl_0_out);

   Delay1No120_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add113_0_impl_0_out,
                 Y => Delay1No120_out);

SharedReg501_out_to_MUX_Add113_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg501_out;
SharedReg21_out_to_MUX_Add113_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg21_out;
SharedReg30_out_to_MUX_Add113_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg30_out;
SharedReg604_out_to_MUX_Add113_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg604_out;
SharedReg939_out_to_MUX_Add113_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg939_out;
SharedReg480_out_to_MUX_Add113_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg480_out;
SharedReg480_out_to_MUX_Add113_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg480_out;
SharedReg158_out_to_MUX_Add113_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg158_out;
SharedReg1004_out_to_MUX_Add113_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1004_out;
SharedReg252_out_to_MUX_Add113_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg252_out;
SharedReg1074_out_to_MUX_Add113_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1074_out;
SharedReg605_out_to_MUX_Add113_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg605_out;
   MUX_Add113_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg501_out_to_MUX_Add113_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg21_out_to_MUX_Add113_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1074_out_to_MUX_Add113_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg605_out_to_MUX_Add113_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg30_out_to_MUX_Add113_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg604_out_to_MUX_Add113_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg939_out_to_MUX_Add113_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg480_out_to_MUX_Add113_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg480_out_to_MUX_Add113_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg158_out_to_MUX_Add113_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1004_out_to_MUX_Add113_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg252_out_to_MUX_Add113_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add113_0_impl_1_out);

   Delay1No121_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add113_0_impl_1_out,
                 Y => Delay1No121_out);

Delay1No122_out_to_Add113_1_impl_parent_implementedSystem_port_0_cast <= Delay1No122_out;
Delay1No123_out_to_Add113_1_impl_parent_implementedSystem_port_1_cast <= Delay1No123_out;
   Add113_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add113_1_impl_out,
                 X => Delay1No122_out_to_Add113_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No123_out_to_Add113_1_impl_parent_implementedSystem_port_1_cast);

SharedReg165_out_to_MUX_Add113_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg165_out;
Delay3No239_out_to_MUX_Add113_1_impl_0_parent_implementedSystem_port_2_cast <= Delay3No239_out;
SharedReg483_out_to_MUX_Add113_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg483_out;
SharedReg5_out_to_MUX_Add113_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg5_out;
SharedReg14_out_to_MUX_Add113_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg14_out;
SharedReg723_out_to_MUX_Add113_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg723_out;
SharedReg553_out_to_MUX_Add113_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg553_out;
SharedReg552_out_to_MUX_Add113_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg552_out;
SharedReg552_out_to_MUX_Add113_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg552_out;
SharedReg418_out_to_MUX_Add113_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg418_out;
SharedReg505_out_to_MUX_Add113_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg505_out;
SharedReg984_out_to_MUX_Add113_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg984_out;
   MUX_Add113_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg165_out_to_MUX_Add113_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay3No239_out_to_MUX_Add113_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg505_out_to_MUX_Add113_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg984_out_to_MUX_Add113_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg483_out_to_MUX_Add113_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg5_out_to_MUX_Add113_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg14_out_to_MUX_Add113_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg723_out_to_MUX_Add113_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg553_out_to_MUX_Add113_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg552_out_to_MUX_Add113_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg552_out_to_MUX_Add113_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg418_out_to_MUX_Add113_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add113_1_impl_0_out);

   Delay1No122_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add113_1_impl_0_out,
                 Y => Delay1No122_out);

SharedReg378_out_to_MUX_Add113_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg378_out;
SharedReg608_out_to_MUX_Add113_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg608_out;
SharedReg505_out_to_MUX_Add113_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg505_out;
SharedReg21_out_to_MUX_Add113_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg21_out;
SharedReg30_out_to_MUX_Add113_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg30_out;
SharedReg804_out_to_MUX_Add113_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg804_out;
SharedReg607_out_to_MUX_Add113_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg607_out;
SharedReg606_out_to_MUX_Add113_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg606_out;
SharedReg606_out_to_MUX_Add113_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg606_out;
SharedReg483_out_to_MUX_Add113_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg483_out;
SharedReg532_out_to_MUX_Add113_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg532_out;
SharedReg443_out_to_MUX_Add113_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg443_out;
   MUX_Add113_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg378_out_to_MUX_Add113_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg608_out_to_MUX_Add113_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg532_out_to_MUX_Add113_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg443_out_to_MUX_Add113_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg505_out_to_MUX_Add113_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg21_out_to_MUX_Add113_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg30_out_to_MUX_Add113_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg804_out_to_MUX_Add113_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg607_out_to_MUX_Add113_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg606_out_to_MUX_Add113_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg606_out_to_MUX_Add113_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg483_out_to_MUX_Add113_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add113_1_impl_1_out);

   Delay1No123_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add113_1_impl_1_out,
                 Y => Delay1No123_out);

Delay1No124_out_to_Add113_2_impl_parent_implementedSystem_port_0_cast <= Delay1No124_out;
Delay1No125_out_to_Add113_2_impl_parent_implementedSystem_port_1_cast <= Delay1No125_out;
   Add113_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add113_2_impl_out,
                 X => Delay1No124_out_to_Add113_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No125_out_to_Add113_2_impl_parent_implementedSystem_port_1_cast);

SharedReg509_out_to_MUX_Add113_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg509_out;
SharedReg260_out_to_MUX_Add113_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg260_out;
SharedReg1013_out_to_MUX_Add113_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1013_out;
SharedReg729_out_to_MUX_Add113_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg729_out;
SharedReg201_out_to_MUX_Add113_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg201_out;
SharedReg5_out_to_MUX_Add113_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg5_out;
SharedReg14_out_to_MUX_Add113_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg14_out;
SharedReg727_out_to_MUX_Add113_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg727_out;
SharedReg555_out_to_MUX_Add113_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg555_out;
SharedReg554_out_to_MUX_Add113_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg554_out;
SharedReg554_out_to_MUX_Add113_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg554_out;
SharedReg420_out_to_MUX_Add113_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg420_out;
   MUX_Add113_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg509_out_to_MUX_Add113_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg260_out_to_MUX_Add113_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg554_out_to_MUX_Add113_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg420_out_to_MUX_Add113_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1013_out_to_MUX_Add113_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg729_out_to_MUX_Add113_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg201_out_to_MUX_Add113_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg5_out_to_MUX_Add113_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg14_out_to_MUX_Add113_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg727_out_to_MUX_Add113_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg555_out_to_MUX_Add113_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg554_out_to_MUX_Add113_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add113_2_impl_0_out);

   Delay1No124_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add113_2_impl_0_out,
                 Y => Delay1No124_out);

SharedReg535_out_to_MUX_Add113_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg535_out;
SharedReg242_out_to_MUX_Add113_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg242_out;
SharedReg1016_out_to_MUX_Add113_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1016_out;
Delay4No184_out_to_MUX_Add113_2_impl_1_parent_implementedSystem_port_4_cast <= Delay4No184_out;
SharedReg349_out_to_MUX_Add113_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg349_out;
SharedReg21_out_to_MUX_Add113_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg21_out;
SharedReg30_out_to_MUX_Add113_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg30_out;
SharedReg807_out_to_MUX_Add113_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg807_out;
SharedReg610_out_to_MUX_Add113_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg610_out;
SharedReg609_out_to_MUX_Add113_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg609_out;
SharedReg609_out_to_MUX_Add113_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg609_out;
SharedReg486_out_to_MUX_Add113_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg486_out;
   MUX_Add113_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg535_out_to_MUX_Add113_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg242_out_to_MUX_Add113_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg609_out_to_MUX_Add113_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg486_out_to_MUX_Add113_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1016_out_to_MUX_Add113_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay4No184_out_to_MUX_Add113_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg349_out_to_MUX_Add113_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg21_out_to_MUX_Add113_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg30_out_to_MUX_Add113_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg807_out_to_MUX_Add113_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg610_out_to_MUX_Add113_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg609_out_to_MUX_Add113_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add113_2_impl_1_out);

   Delay1No125_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add113_2_impl_1_out,
                 Y => Delay1No125_out);

Delay1No126_out_to_Add113_3_impl_parent_implementedSystem_port_0_cast <= Delay1No126_out;
Delay1No127_out_to_Add113_3_impl_parent_implementedSystem_port_1_cast <= Delay1No127_out;
   Add113_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add113_3_impl_out,
                 X => Delay1No126_out_to_Add113_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No127_out_to_Add113_3_impl_parent_implementedSystem_port_1_cast);

SharedReg556_out_to_MUX_Add113_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg556_out;
SharedReg513_out_to_MUX_Add113_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg513_out;
SharedReg861_out_to_MUX_Add113_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg861_out;
SharedReg1018_out_to_MUX_Add113_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1018_out;
Delay3No241_out_to_MUX_Add113_3_impl_0_parent_implementedSystem_port_5_cast <= Delay3No241_out;
SharedReg489_out_to_MUX_Add113_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg489_out;
SharedReg5_out_to_MUX_Add113_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg5_out;
SharedReg405_out_to_MUX_Add113_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg405_out;
SharedReg731_out_to_MUX_Add113_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg731_out;
SharedReg731_out_to_MUX_Add113_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg731_out;
SharedReg730_out_to_MUX_Add113_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg730_out;
SharedReg730_out_to_MUX_Add113_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg730_out;
   MUX_Add113_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg556_out_to_MUX_Add113_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg513_out_to_MUX_Add113_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg730_out_to_MUX_Add113_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg730_out_to_MUX_Add113_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg861_out_to_MUX_Add113_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1018_out_to_MUX_Add113_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay3No241_out_to_MUX_Add113_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg489_out_to_MUX_Add113_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg5_out_to_MUX_Add113_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg405_out_to_MUX_Add113_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg731_out_to_MUX_Add113_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg731_out_to_MUX_Add113_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add113_3_impl_0_out);

   Delay1No126_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add113_3_impl_0_out,
                 Y => Delay1No126_out);

SharedReg612_out_to_MUX_Add113_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg612_out;
SharedReg538_out_to_MUX_Add113_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg538_out;
SharedReg756_out_to_MUX_Add113_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg756_out;
SharedReg1021_out_to_MUX_Add113_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1021_out;
SharedReg614_out_to_MUX_Add113_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg614_out;
SharedReg513_out_to_MUX_Add113_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg513_out;
SharedReg21_out_to_MUX_Add113_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg21_out;
SharedReg733_out_to_MUX_Add113_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg733_out;
SharedReg810_out_to_MUX_Add113_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg810_out;
SharedReg810_out_to_MUX_Add113_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg810_out;
SharedReg809_out_to_MUX_Add113_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg809_out;
SharedReg809_out_to_MUX_Add113_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg809_out;
   MUX_Add113_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg612_out_to_MUX_Add113_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg538_out_to_MUX_Add113_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg809_out_to_MUX_Add113_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg809_out_to_MUX_Add113_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg756_out_to_MUX_Add113_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1021_out_to_MUX_Add113_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg614_out_to_MUX_Add113_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg513_out_to_MUX_Add113_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg21_out_to_MUX_Add113_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg733_out_to_MUX_Add113_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg810_out_to_MUX_Add113_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg810_out_to_MUX_Add113_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add113_3_impl_1_out);

   Delay1No127_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add113_3_impl_1_out,
                 Y => Delay1No127_out);

Delay1No128_out_to_Add113_4_impl_parent_implementedSystem_port_0_cast <= Delay1No128_out;
Delay1No129_out_to_Add113_4_impl_parent_implementedSystem_port_1_cast <= Delay1No129_out;
   Add113_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add113_4_impl_out,
                 X => Delay1No128_out_to_Add113_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No129_out_to_Add113_4_impl_parent_implementedSystem_port_1_cast);

SharedReg734_out_to_MUX_Add113_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg734_out;
SharedReg558_out_to_MUX_Add113_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg558_out;
SharedReg424_out_to_MUX_Add113_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg424_out;
SharedReg461_out_to_MUX_Add113_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg461_out;
SharedReg206_out_to_MUX_Add113_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg206_out;
SharedReg994_out_to_MUX_Add113_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg994_out;
SharedReg737_out_to_MUX_Add113_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg737_out;
SharedReg492_out_to_MUX_Add113_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg492_out;
SharedReg5_out_to_MUX_Add113_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg5_out;
SharedReg408_out_to_MUX_Add113_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg408_out;
SharedReg928_out_to_MUX_Add113_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg928_out;
SharedReg735_out_to_MUX_Add113_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg735_out;
   MUX_Add113_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg734_out_to_MUX_Add113_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg558_out_to_MUX_Add113_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg928_out_to_MUX_Add113_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg735_out_to_MUX_Add113_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg424_out_to_MUX_Add113_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg461_out_to_MUX_Add113_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg206_out_to_MUX_Add113_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg994_out_to_MUX_Add113_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg737_out_to_MUX_Add113_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg492_out_to_MUX_Add113_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg5_out_to_MUX_Add113_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg408_out_to_MUX_Add113_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add113_4_impl_0_out);

   Delay1No128_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add113_4_impl_0_out,
                 Y => Delay1No128_out);

SharedReg812_out_to_MUX_Add113_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg812_out;
SharedReg615_out_to_MUX_Add113_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg615_out;
SharedReg492_out_to_MUX_Add113_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg492_out;
SharedReg689_out_to_MUX_Add113_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg689_out;
SharedReg211_out_to_MUX_Add113_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg211_out;
SharedReg1027_out_to_MUX_Add113_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1027_out;
Delay4No186_out_to_MUX_Add113_4_impl_1_parent_implementedSystem_port_7_cast <= Delay4No186_out;
SharedReg517_out_to_MUX_Add113_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg517_out;
SharedReg21_out_to_MUX_Add113_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg21_out;
SharedReg737_out_to_MUX_Add113_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg737_out;
SharedReg952_out_to_MUX_Add113_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg952_out;
SharedReg813_out_to_MUX_Add113_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg813_out;
   MUX_Add113_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg812_out_to_MUX_Add113_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg615_out_to_MUX_Add113_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg952_out_to_MUX_Add113_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg813_out_to_MUX_Add113_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg492_out_to_MUX_Add113_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg689_out_to_MUX_Add113_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg211_out_to_MUX_Add113_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1027_out_to_MUX_Add113_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay4No186_out_to_MUX_Add113_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg517_out_to_MUX_Add113_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg21_out_to_MUX_Add113_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg737_out_to_MUX_Add113_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add113_4_impl_1_out);

   Delay1No129_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add113_4_impl_1_out,
                 Y => Delay1No129_out);

Delay1No130_out_to_Add24_5_impl_parent_implementedSystem_port_0_cast <= Delay1No130_out;
Delay1No131_out_to_Add24_5_impl_parent_implementedSystem_port_1_cast <= Delay1No131_out;
   Add24_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add24_5_impl_out,
                 X => Delay1No130_out_to_Add24_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No131_out_to_Add24_5_impl_parent_implementedSystem_port_1_cast);

SharedReg769_out_to_MUX_Add24_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg769_out;
SharedReg927_out_to_MUX_Add24_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg927_out;
SharedReg734_out_to_MUX_Add24_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg734_out;
SharedReg927_out_to_MUX_Add24_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg927_out;
SharedReg272_out_to_MUX_Add24_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg272_out;
SharedReg657_out_to_MUX_Add24_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg657_out;
SharedReg736_out_to_MUX_Add24_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg736_out;
Delay4No221_out_to_MUX_Add24_5_impl_0_parent_implementedSystem_port_8_cast <= Delay4No221_out;
SharedReg10_out_to_MUX_Add24_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg10_out;
SharedReg839_out_to_MUX_Add24_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg839_out;
SharedReg974_out_to_MUX_Add24_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg974_out;
SharedReg928_out_to_MUX_Add24_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg928_out;
   MUX_Add24_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg769_out_to_MUX_Add24_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg927_out_to_MUX_Add24_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg974_out_to_MUX_Add24_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg928_out_to_MUX_Add24_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg734_out_to_MUX_Add24_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg927_out_to_MUX_Add24_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg272_out_to_MUX_Add24_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg657_out_to_MUX_Add24_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg736_out_to_MUX_Add24_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay4No221_out_to_MUX_Add24_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg10_out_to_MUX_Add24_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg839_out_to_MUX_Add24_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add24_5_impl_0_out);

   Delay1No130_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add24_5_impl_0_out,
                 Y => Delay1No130_out);

SharedReg714_out_to_MUX_Add24_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg714_out;
SharedReg951_out_to_MUX_Add24_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg951_out;
SharedReg812_out_to_MUX_Add24_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg812_out;
SharedReg951_out_to_MUX_Add24_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg951_out;
SharedReg276_out_to_MUX_Add24_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg276_out;
SharedReg734_out_to_MUX_Add24_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg734_out;
SharedReg814_out_to_MUX_Add24_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg814_out;
Delay4No228_out_to_MUX_Add24_5_impl_1_parent_implementedSystem_port_8_cast <= Delay4No228_out;
SharedReg26_out_to_MUX_Add24_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg26_out;
SharedReg637_out_to_MUX_Add24_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg637_out;
SharedReg930_out_to_MUX_Add24_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg930_out;
SharedReg952_out_to_MUX_Add24_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg952_out;
   MUX_Add24_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg714_out_to_MUX_Add24_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg951_out_to_MUX_Add24_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg930_out_to_MUX_Add24_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg952_out_to_MUX_Add24_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg812_out_to_MUX_Add24_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg951_out_to_MUX_Add24_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg276_out_to_MUX_Add24_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg734_out_to_MUX_Add24_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg814_out_to_MUX_Add24_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay4No228_out_to_MUX_Add24_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg26_out_to_MUX_Add24_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg637_out_to_MUX_Add24_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add24_5_impl_1_out);

   Delay1No131_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add24_5_impl_1_out,
                 Y => Delay1No131_out);

Delay1No132_out_to_Add32_5_impl_parent_implementedSystem_port_0_cast <= Delay1No132_out;
Delay1No133_out_to_Add32_5_impl_parent_implementedSystem_port_1_cast <= Delay1No133_out;
   Add32_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add32_5_impl_out,
                 X => Delay1No132_out_to_Add32_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No133_out_to_Add32_5_impl_parent_implementedSystem_port_1_cast);

SharedReg932_out_to_MUX_Add32_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg932_out;
SharedReg561_out_to_MUX_Add32_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg561_out;
SharedReg560_out_to_MUX_Add32_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg560_out;
SharedReg426_out_to_MUX_Add32_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg426_out;
SharedReg152_out_to_MUX_Add32_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg152_out;
SharedReg468_out_to_MUX_Add32_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg468_out;
SharedReg694_out_to_MUX_Add32_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg694_out;
SharedReg1029_out_to_MUX_Add32_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1029_out;
SharedReg741_out_to_MUX_Add32_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg741_out;
SharedReg495_out_to_MUX_Add32_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg495_out;
SharedReg6_out_to_MUX_Add32_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg6_out;
SharedReg411_out_to_MUX_Add32_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg411_out;
   MUX_Add32_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg932_out_to_MUX_Add32_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg561_out_to_MUX_Add32_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg6_out_to_MUX_Add32_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg411_out_to_MUX_Add32_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg560_out_to_MUX_Add32_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg426_out_to_MUX_Add32_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg152_out_to_MUX_Add32_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg468_out_to_MUX_Add32_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg694_out_to_MUX_Add32_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1029_out_to_MUX_Add32_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg741_out_to_MUX_Add32_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg495_out_to_MUX_Add32_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add32_5_impl_0_out);

   Delay1No132_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add32_5_impl_0_out,
                 Y => Delay1No132_out);

SharedReg955_out_to_MUX_Add32_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg955_out;
SharedReg619_out_to_MUX_Add32_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg619_out;
SharedReg618_out_to_MUX_Add32_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg618_out;
SharedReg495_out_to_MUX_Add32_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg495_out;
SharedReg224_out_to_MUX_Add32_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg224_out;
SharedReg694_out_to_MUX_Add32_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg694_out;
SharedReg716_out_to_MUX_Add32_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg716_out;
SharedReg1065_out_to_MUX_Add32_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1065_out;
Delay4No187_out_to_MUX_Add32_5_impl_1_parent_implementedSystem_port_9_cast <= Delay4No187_out;
SharedReg521_out_to_MUX_Add32_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg521_out;
SharedReg22_out_to_MUX_Add32_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg22_out;
SharedReg741_out_to_MUX_Add32_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg741_out;
   MUX_Add32_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg955_out_to_MUX_Add32_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg619_out_to_MUX_Add32_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg22_out_to_MUX_Add32_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg741_out_to_MUX_Add32_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg618_out_to_MUX_Add32_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg495_out_to_MUX_Add32_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg224_out_to_MUX_Add32_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg694_out_to_MUX_Add32_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg716_out_to_MUX_Add32_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1065_out_to_MUX_Add32_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay4No187_out_to_MUX_Add32_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg521_out_to_MUX_Add32_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add32_5_impl_1_out);

   Delay1No133_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add32_5_impl_1_out,
                 Y => Delay1No133_out);

Delay1No134_out_to_Add122_5_impl_parent_implementedSystem_port_0_cast <= Delay1No134_out;
Delay1No135_out_to_Add122_5_impl_parent_implementedSystem_port_1_cast <= Delay1No135_out;
   Add122_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add122_5_impl_out,
                 X => Delay1No134_out_to_Add122_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No135_out_to_Add122_5_impl_parent_implementedSystem_port_1_cast);

Delay6No47_out_to_MUX_Add122_5_impl_0_parent_implementedSystem_port_1_cast <= Delay6No47_out;
SharedReg739_out_to_MUX_Add122_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg739_out;
SharedReg738_out_to_MUX_Add122_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg738_out;
SharedReg560_out_to_MUX_Add122_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg560_out;
SharedReg426_out_to_MUX_Add122_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg426_out;
SharedReg521_out_to_MUX_Add122_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg521_out;
SharedReg286_out_to_MUX_Add122_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg286_out;
SharedReg225_out_to_MUX_Add122_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg225_out;
Delay3No243_out_to_MUX_Add122_5_impl_0_parent_implementedSystem_port_9_cast <= Delay3No243_out;
SharedReg560_out_to_MUX_Add122_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg560_out;
SharedReg10_out_to_MUX_Add122_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg10_out;
SharedReg545_out_to_MUX_Add122_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg545_out;
   MUX_Add122_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay6No47_out_to_MUX_Add122_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg739_out_to_MUX_Add122_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg10_out_to_MUX_Add122_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg545_out_to_MUX_Add122_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg738_out_to_MUX_Add122_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg560_out_to_MUX_Add122_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg426_out_to_MUX_Add122_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg521_out_to_MUX_Add122_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg286_out_to_MUX_Add122_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg225_out_to_MUX_Add122_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay3No243_out_to_MUX_Add122_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg560_out_to_MUX_Add122_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add122_5_impl_0_out);

   Delay1No134_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add122_5_impl_0_out,
                 Y => Delay1No134_out);

SharedReg933_out_to_MUX_Add122_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg933_out;
SharedReg816_out_to_MUX_Add122_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg816_out;
SharedReg815_out_to_MUX_Add122_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg815_out;
SharedReg618_out_to_MUX_Add122_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg618_out;
SharedReg495_out_to_MUX_Add122_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg495_out;
SharedReg544_out_to_MUX_Add122_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg544_out;
SharedReg289_out_to_MUX_Add122_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg289_out;
SharedReg231_out_to_MUX_Add122_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg231_out;
SharedReg620_out_to_MUX_Add122_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg620_out;
SharedReg618_out_to_MUX_Add122_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg618_out;
SharedReg26_out_to_MUX_Add122_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg26_out;
SharedReg817_out_to_MUX_Add122_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg817_out;
   MUX_Add122_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg933_out_to_MUX_Add122_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg816_out_to_MUX_Add122_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg26_out_to_MUX_Add122_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg817_out_to_MUX_Add122_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg815_out_to_MUX_Add122_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg618_out_to_MUX_Add122_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg495_out_to_MUX_Add122_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg544_out_to_MUX_Add122_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg289_out_to_MUX_Add122_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg231_out_to_MUX_Add122_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg620_out_to_MUX_Add122_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg618_out_to_MUX_Add122_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add122_5_impl_1_out);

   Delay1No135_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add122_5_impl_1_out,
                 Y => Delay1No135_out);

Delay1No136_out_to_Add33_0_impl_parent_implementedSystem_port_0_cast <= Delay1No136_out;
Delay1No137_out_to_Add33_0_impl_parent_implementedSystem_port_1_cast <= Delay1No137_out;
   Add33_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add33_0_impl_out,
                 X => Delay1No136_out_to_Add33_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No137_out_to_Add33_0_impl_parent_implementedSystem_port_1_cast);

SharedReg550_out_to_MUX_Add33_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg550_out;
SharedReg6_out_to_MUX_Add33_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg6_out;
SharedReg396_out_to_MUX_Add33_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg396_out;
SharedReg719_out_to_MUX_Add33_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg719_out;
SharedReg551_out_to_MUX_Add33_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg551_out;
SharedReg550_out_to_MUX_Add33_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg550_out;
SharedReg550_out_to_MUX_Add33_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg550_out;
SharedReg416_out_to_MUX_Add33_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg416_out;
SharedReg501_out_to_MUX_Add33_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg501_out;
SharedReg1004_out_to_MUX_Add33_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1004_out;
SharedReg159_out_to_MUX_Add33_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg159_out;
SharedReg720_out_to_MUX_Add33_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg720_out;
   MUX_Add33_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg550_out_to_MUX_Add33_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg6_out_to_MUX_Add33_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg159_out_to_MUX_Add33_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg720_out_to_MUX_Add33_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg396_out_to_MUX_Add33_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg719_out_to_MUX_Add33_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg551_out_to_MUX_Add33_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg550_out_to_MUX_Add33_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg550_out_to_MUX_Add33_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg416_out_to_MUX_Add33_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg501_out_to_MUX_Add33_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1004_out_to_MUX_Add33_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add33_0_impl_0_out);

   Delay1No136_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add33_0_impl_0_out,
                 Y => Delay1No136_out);

SharedReg603_out_to_MUX_Add33_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg603_out;
SharedReg22_out_to_MUX_Add33_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg22_out;
SharedReg721_out_to_MUX_Add33_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg721_out;
SharedReg801_out_to_MUX_Add33_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg801_out;
SharedReg604_out_to_MUX_Add33_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg604_out;
SharedReg603_out_to_MUX_Add33_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg603_out;
SharedReg603_out_to_MUX_Add33_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg603_out;
SharedReg480_out_to_MUX_Add33_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg480_out;
SharedReg529_out_to_MUX_Add33_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg529_out;
SharedReg568_out_to_MUX_Add33_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg568_out;
SharedReg369_out_to_MUX_Add33_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg369_out;
SharedReg802_out_to_MUX_Add33_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg802_out;
   MUX_Add33_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg603_out_to_MUX_Add33_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg22_out_to_MUX_Add33_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg369_out_to_MUX_Add33_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg802_out_to_MUX_Add33_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg721_out_to_MUX_Add33_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg801_out_to_MUX_Add33_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg604_out_to_MUX_Add33_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg603_out_to_MUX_Add33_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg603_out_to_MUX_Add33_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg480_out_to_MUX_Add33_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg529_out_to_MUX_Add33_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg568_out_to_MUX_Add33_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add33_0_impl_1_out);

   Delay1No137_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add33_0_impl_1_out,
                 Y => Delay1No137_out);

Delay1No138_out_to_Add33_2_impl_parent_implementedSystem_port_0_cast <= Delay1No138_out;
Delay1No139_out_to_Add33_2_impl_parent_implementedSystem_port_1_cast <= Delay1No139_out;
   Add33_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add33_2_impl_out,
                 X => Delay1No138_out_to_Add33_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No139_out_to_Add33_2_impl_parent_implementedSystem_port_1_cast);

SharedReg919_out_to_MUX_Add33_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg919_out;
SharedReg858_out_to_MUX_Add33_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg858_out;
SharedReg171_out_to_MUX_Add33_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg171_out;
Delay3No240_out_to_MUX_Add33_2_impl_0_parent_implementedSystem_port_4_cast <= Delay3No240_out;
SharedReg486_out_to_MUX_Add33_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg486_out;
SharedReg6_out_to_MUX_Add33_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg6_out;
SharedReg402_out_to_MUX_Add33_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg402_out;
SharedReg920_out_to_MUX_Add33_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg920_out;
SharedReg727_out_to_MUX_Add33_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg727_out;
SharedReg726_out_to_MUX_Add33_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg726_out;
SharedReg726_out_to_MUX_Add33_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg726_out;
SharedReg554_out_to_MUX_Add33_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg554_out;
   MUX_Add33_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg919_out_to_MUX_Add33_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg858_out_to_MUX_Add33_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg726_out_to_MUX_Add33_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg554_out_to_MUX_Add33_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg171_out_to_MUX_Add33_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay3No240_out_to_MUX_Add33_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg486_out_to_MUX_Add33_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg6_out_to_MUX_Add33_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg402_out_to_MUX_Add33_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg920_out_to_MUX_Add33_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg727_out_to_MUX_Add33_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg726_out_to_MUX_Add33_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add33_2_impl_0_out);

   Delay1No138_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add33_2_impl_0_out,
                 Y => Delay1No138_out);

SharedReg945_out_to_MUX_Add33_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg945_out;
SharedReg751_out_to_MUX_Add33_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg751_out;
SharedReg347_out_to_MUX_Add33_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg347_out;
SharedReg611_out_to_MUX_Add33_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg611_out;
SharedReg509_out_to_MUX_Add33_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg509_out;
SharedReg22_out_to_MUX_Add33_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg22_out;
SharedReg729_out_to_MUX_Add33_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg729_out;
SharedReg946_out_to_MUX_Add33_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg946_out;
SharedReg807_out_to_MUX_Add33_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg807_out;
SharedReg806_out_to_MUX_Add33_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg806_out;
SharedReg806_out_to_MUX_Add33_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg806_out;
SharedReg609_out_to_MUX_Add33_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg609_out;
   MUX_Add33_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg945_out_to_MUX_Add33_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg751_out_to_MUX_Add33_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg806_out_to_MUX_Add33_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg609_out_to_MUX_Add33_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg347_out_to_MUX_Add33_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg611_out_to_MUX_Add33_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg509_out_to_MUX_Add33_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg22_out_to_MUX_Add33_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg729_out_to_MUX_Add33_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg946_out_to_MUX_Add33_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg807_out_to_MUX_Add33_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg806_out_to_MUX_Add33_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add33_2_impl_1_out);

   Delay1No139_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add33_2_impl_1_out,
                 Y => Delay1No139_out);

Delay1No140_out_to_Add33_4_impl_parent_implementedSystem_port_0_cast <= Delay1No140_out;
Delay1No141_out_to_Add33_4_impl_parent_implementedSystem_port_1_cast <= Delay1No141_out;
   Add33_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add33_4_impl_out,
                 X => Delay1No140_out_to_Add33_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No141_out_to_Add33_4_impl_parent_implementedSystem_port_1_cast);

SharedReg927_out_to_MUX_Add33_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg927_out;
SharedReg734_out_to_MUX_Add33_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg734_out;
SharedReg558_out_to_MUX_Add33_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg558_out;
SharedReg517_out_to_MUX_Add33_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg517_out;
SharedReg689_out_to_MUX_Add33_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg689_out;
SharedReg279_out_to_MUX_Add33_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg279_out;
Delay3No242_out_to_MUX_Add33_4_impl_0_parent_implementedSystem_port_7_cast <= Delay3No242_out;
SharedReg558_out_to_MUX_Add33_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg558_out;
SharedReg6_out_to_MUX_Add33_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg6_out;
SharedReg542_out_to_MUX_Add33_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg542_out;
Delay6No46_out_to_MUX_Add33_4_impl_0_parent_implementedSystem_port_11_cast <= Delay6No46_out;
SharedReg425_out_to_MUX_Add33_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg425_out;
   MUX_Add33_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg927_out_to_MUX_Add33_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg734_out_to_MUX_Add33_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay6No46_out_to_MUX_Add33_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg425_out_to_MUX_Add33_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg558_out_to_MUX_Add33_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg517_out_to_MUX_Add33_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg689_out_to_MUX_Add33_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg279_out_to_MUX_Add33_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay3No242_out_to_MUX_Add33_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg558_out_to_MUX_Add33_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg6_out_to_MUX_Add33_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg542_out_to_MUX_Add33_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add33_4_impl_0_out);

   Delay1No140_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add33_4_impl_0_out,
                 Y => Delay1No140_out);

SharedReg951_out_to_MUX_Add33_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg951_out;
SharedReg812_out_to_MUX_Add33_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg812_out;
SharedReg615_out_to_MUX_Add33_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg615_out;
SharedReg541_out_to_MUX_Add33_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg541_out;
SharedReg710_out_to_MUX_Add33_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg710_out;
SharedReg284_out_to_MUX_Add33_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg284_out;
SharedReg617_out_to_MUX_Add33_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg617_out;
SharedReg615_out_to_MUX_Add33_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg615_out;
SharedReg22_out_to_MUX_Add33_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg22_out;
SharedReg814_out_to_MUX_Add33_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg814_out;
SharedReg929_out_to_MUX_Add33_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg929_out;
SharedReg493_out_to_MUX_Add33_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg493_out;
   MUX_Add33_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg951_out_to_MUX_Add33_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg812_out_to_MUX_Add33_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg929_out_to_MUX_Add33_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg493_out_to_MUX_Add33_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg615_out_to_MUX_Add33_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg541_out_to_MUX_Add33_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg710_out_to_MUX_Add33_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg284_out_to_MUX_Add33_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg617_out_to_MUX_Add33_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg615_out_to_MUX_Add33_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg22_out_to_MUX_Add33_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg814_out_to_MUX_Add33_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add33_4_impl_1_out);

   Delay1No141_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add33_4_impl_1_out,
                 Y => Delay1No141_out);

Delay1No142_out_to_Add33_5_impl_parent_implementedSystem_port_0_cast <= Delay1No142_out;
Delay1No143_out_to_Add33_5_impl_parent_implementedSystem_port_1_cast <= Delay1No143_out;
   Add33_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add33_5_impl_out,
                 X => Delay1No142_out_to_Add33_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No143_out_to_Add33_5_impl_parent_implementedSystem_port_1_cast);

SharedReg977_out_to_MUX_Add33_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg977_out;
SharedReg427_out_to_MUX_Add33_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg427_out;
SharedReg931_out_to_MUX_Add33_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg931_out;
SharedReg738_out_to_MUX_Add33_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg738_out;
SharedReg560_out_to_MUX_Add33_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg560_out;
SharedReg931_out_to_MUX_Add33_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg931_out;
SharedReg868_out_to_MUX_Add33_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg868_out;
SharedReg660_out_to_MUX_Add33_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg660_out;
SharedReg740_out_to_MUX_Add33_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg740_out;
Delay4No222_out_to_MUX_Add33_5_impl_0_parent_implementedSystem_port_10_cast <= Delay4No222_out;
SharedReg13_out_to_MUX_Add33_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg13_out;
SharedReg843_out_to_MUX_Add33_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg843_out;
   MUX_Add33_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg977_out_to_MUX_Add33_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg427_out_to_MUX_Add33_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg13_out_to_MUX_Add33_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg843_out_to_MUX_Add33_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg931_out_to_MUX_Add33_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg738_out_to_MUX_Add33_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg560_out_to_MUX_Add33_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg931_out_to_MUX_Add33_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg868_out_to_MUX_Add33_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg660_out_to_MUX_Add33_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg740_out_to_MUX_Add33_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay4No222_out_to_MUX_Add33_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add33_5_impl_0_out);

   Delay1No142_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add33_5_impl_0_out,
                 Y => Delay1No142_out);

SharedReg934_out_to_MUX_Add33_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg934_out;
SharedReg496_out_to_MUX_Add33_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg496_out;
SharedReg954_out_to_MUX_Add33_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg954_out;
SharedReg815_out_to_MUX_Add33_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg815_out;
SharedReg618_out_to_MUX_Add33_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg618_out;
SharedReg954_out_to_MUX_Add33_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg954_out;
SharedReg471_out_to_MUX_Add33_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg471_out;
SharedReg738_out_to_MUX_Add33_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg738_out;
SharedReg817_out_to_MUX_Add33_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg817_out;
Delay4No229_out_to_MUX_Add33_5_impl_1_parent_implementedSystem_port_10_cast <= Delay4No229_out;
SharedReg29_out_to_MUX_Add33_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg29_out;
SharedReg640_out_to_MUX_Add33_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg640_out;
   MUX_Add33_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg934_out_to_MUX_Add33_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg496_out_to_MUX_Add33_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg29_out_to_MUX_Add33_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg640_out_to_MUX_Add33_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg954_out_to_MUX_Add33_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg815_out_to_MUX_Add33_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg618_out_to_MUX_Add33_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg954_out_to_MUX_Add33_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg471_out_to_MUX_Add33_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg738_out_to_MUX_Add33_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg817_out_to_MUX_Add33_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay4No229_out_to_MUX_Add33_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add33_5_impl_1_out);

   Delay1No143_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add33_5_impl_1_out,
                 Y => Delay1No143_out);

Delay1No144_out_to_Add33_6_impl_parent_implementedSystem_port_0_cast <= Delay1No144_out;
Delay1No145_out_to_Add33_6_impl_parent_implementedSystem_port_1_cast <= Delay1No145_out;
   Add33_6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add33_6_impl_out,
                 X => Delay1No144_out_to_Add33_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No145_out_to_Add33_6_impl_parent_implementedSystem_port_1_cast);

SharedReg548_out_to_MUX_Add33_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg548_out;
SharedReg743_out_to_MUX_Add33_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg743_out;
SharedReg743_out_to_MUX_Add33_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg743_out;
SharedReg562_out_to_MUX_Add33_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg562_out;
SharedReg562_out_to_MUX_Add33_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg562_out;
SharedReg428_out_to_MUX_Add33_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg428_out;
SharedReg476_out_to_MUX_Add33_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg476_out;
SharedReg1001_out_to_MUX_Add33_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1001_out;
SharedReg1067_out_to_MUX_Add33_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1067_out;
SharedReg744_out_to_MUX_Add33_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg744_out;
SharedReg562_out_to_MUX_Add33_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg562_out;
SharedReg6_out_to_MUX_Add33_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg6_out;
   MUX_Add33_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg548_out_to_MUX_Add33_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg743_out_to_MUX_Add33_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg562_out_to_MUX_Add33_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg6_out_to_MUX_Add33_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg743_out_to_MUX_Add33_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg562_out_to_MUX_Add33_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg562_out_to_MUX_Add33_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg428_out_to_MUX_Add33_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg476_out_to_MUX_Add33_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1001_out_to_MUX_Add33_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1067_out_to_MUX_Add33_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg744_out_to_MUX_Add33_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add33_6_impl_0_out);

   Delay1No144_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add33_6_impl_0_out,
                 Y => Delay1No144_out);

SharedReg820_out_to_MUX_Add33_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg820_out;
SharedReg819_out_to_MUX_Add33_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg819_out;
SharedReg819_out_to_MUX_Add33_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg819_out;
SharedReg621_out_to_MUX_Add33_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg621_out;
SharedReg621_out_to_MUX_Add33_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg621_out;
SharedReg498_out_to_MUX_Add33_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg498_out;
SharedReg1033_out_to_MUX_Add33_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1033_out;
SharedReg601_out_to_MUX_Add33_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg601_out;
SharedReg1080_out_to_MUX_Add33_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1080_out;
SharedReg820_out_to_MUX_Add33_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg820_out;
SharedReg621_out_to_MUX_Add33_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg621_out;
SharedReg22_out_to_MUX_Add33_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg22_out;
   MUX_Add33_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg820_out_to_MUX_Add33_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg819_out_to_MUX_Add33_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg621_out_to_MUX_Add33_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg22_out_to_MUX_Add33_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg819_out_to_MUX_Add33_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg621_out_to_MUX_Add33_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg621_out_to_MUX_Add33_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg498_out_to_MUX_Add33_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1033_out_to_MUX_Add33_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg601_out_to_MUX_Add33_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1080_out_to_MUX_Add33_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg820_out_to_MUX_Add33_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add33_6_impl_1_out);

   Delay1No145_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add33_6_impl_1_out,
                 Y => Delay1No145_out);

Delay1No146_out_to_Add123_0_impl_parent_implementedSystem_port_0_cast <= Delay1No146_out;
Delay1No147_out_to_Add123_0_impl_parent_implementedSystem_port_1_cast <= Delay1No147_out;
   Add123_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add123_0_impl_out,
                 X => Delay1No146_out_to_Add123_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No147_out_to_Add123_0_impl_parent_implementedSystem_port_1_cast);

Delay4No217_out_to_MUX_Add123_0_impl_0_parent_implementedSystem_port_1_cast <= Delay4No217_out;
SharedReg10_out_to_MUX_Add123_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg10_out;
SharedReg530_out_to_MUX_Add123_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg530_out;
SharedReg912_out_to_MUX_Add123_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg912_out;
SharedReg719_out_to_MUX_Add123_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg719_out;
SharedReg718_out_to_MUX_Add123_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg718_out;
SharedReg718_out_to_MUX_Add123_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg718_out;
SharedReg550_out_to_MUX_Add123_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg550_out;
SharedReg911_out_to_MUX_Add123_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg911_out;
SharedReg326_out_to_MUX_Add123_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg326_out;
SharedReg645_out_to_MUX_Add123_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg645_out;
SharedReg911_out_to_MUX_Add123_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg911_out;
   MUX_Add123_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay4No217_out_to_MUX_Add123_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg10_out_to_MUX_Add123_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg645_out_to_MUX_Add123_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg911_out_to_MUX_Add123_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg530_out_to_MUX_Add123_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg912_out_to_MUX_Add123_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg719_out_to_MUX_Add123_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg718_out_to_MUX_Add123_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg718_out_to_MUX_Add123_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg550_out_to_MUX_Add123_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg911_out_to_MUX_Add123_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg326_out_to_MUX_Add123_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add123_0_impl_0_out);

   Delay1No146_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add123_0_impl_0_out,
                 Y => Delay1No146_out);

Delay4No224_out_to_MUX_Add123_0_impl_1_parent_implementedSystem_port_1_cast <= Delay4No224_out;
SharedReg26_out_to_MUX_Add123_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg26_out;
SharedReg802_out_to_MUX_Add123_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg802_out;
SharedReg940_out_to_MUX_Add123_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg940_out;
SharedReg801_out_to_MUX_Add123_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg801_out;
SharedReg800_out_to_MUX_Add123_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg800_out;
SharedReg800_out_to_MUX_Add123_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg800_out;
SharedReg603_out_to_MUX_Add123_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg603_out;
SharedReg939_out_to_MUX_Add123_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg939_out;
SharedReg300_out_to_MUX_Add123_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg300_out;
SharedReg718_out_to_MUX_Add123_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg718_out;
SharedReg884_out_to_MUX_Add123_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg884_out;
   MUX_Add123_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay4No224_out_to_MUX_Add123_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg26_out_to_MUX_Add123_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg718_out_to_MUX_Add123_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg884_out_to_MUX_Add123_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg802_out_to_MUX_Add123_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg940_out_to_MUX_Add123_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg801_out_to_MUX_Add123_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg800_out_to_MUX_Add123_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg800_out_to_MUX_Add123_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg603_out_to_MUX_Add123_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg939_out_to_MUX_Add123_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg300_out_to_MUX_Add123_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add123_0_impl_1_out);

   Delay1No147_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add123_0_impl_1_out,
                 Y => Delay1No147_out);

Delay1No148_out_to_Add123_1_impl_parent_implementedSystem_port_0_cast <= Delay1No148_out;
Delay1No149_out_to_Add123_1_impl_parent_implementedSystem_port_1_cast <= Delay1No149_out;
   Add123_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add123_1_impl_out,
                 X => Delay1No148_out_to_Add123_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No149_out_to_Add123_1_impl_parent_implementedSystem_port_1_cast);

SharedReg648_out_to_MUX_Add123_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg648_out;
SharedReg724_out_to_MUX_Add123_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg724_out;
SharedReg552_out_to_MUX_Add123_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg552_out;
SharedReg6_out_to_MUX_Add123_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg6_out;
SharedReg399_out_to_MUX_Add123_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg399_out;
SharedReg916_out_to_MUX_Add123_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg916_out;
SharedReg723_out_to_MUX_Add123_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg723_out;
SharedReg722_out_to_MUX_Add123_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg722_out;
SharedReg722_out_to_MUX_Add123_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg722_out;
SharedReg552_out_to_MUX_Add123_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg552_out;
SharedReg915_out_to_MUX_Add123_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg915_out;
SharedReg335_out_to_MUX_Add123_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg335_out;
   MUX_Add123_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg648_out_to_MUX_Add123_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg724_out_to_MUX_Add123_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg915_out_to_MUX_Add123_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg335_out_to_MUX_Add123_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg552_out_to_MUX_Add123_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg6_out_to_MUX_Add123_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg399_out_to_MUX_Add123_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg916_out_to_MUX_Add123_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg723_out_to_MUX_Add123_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg722_out_to_MUX_Add123_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg722_out_to_MUX_Add123_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg552_out_to_MUX_Add123_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add123_1_impl_0_out);

   Delay1No148_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add123_1_impl_0_out,
                 Y => Delay1No148_out);

SharedReg722_out_to_MUX_Add123_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg722_out;
SharedReg805_out_to_MUX_Add123_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg805_out;
SharedReg606_out_to_MUX_Add123_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg606_out;
SharedReg22_out_to_MUX_Add123_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg22_out;
SharedReg725_out_to_MUX_Add123_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg725_out;
SharedReg943_out_to_MUX_Add123_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg943_out;
SharedReg804_out_to_MUX_Add123_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg804_out;
SharedReg803_out_to_MUX_Add123_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg803_out;
SharedReg803_out_to_MUX_Add123_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg803_out;
SharedReg606_out_to_MUX_Add123_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg606_out;
SharedReg942_out_to_MUX_Add123_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg942_out;
SharedReg258_out_to_MUX_Add123_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg258_out;
   MUX_Add123_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg722_out_to_MUX_Add123_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg805_out_to_MUX_Add123_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg942_out_to_MUX_Add123_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg258_out_to_MUX_Add123_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg606_out_to_MUX_Add123_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg22_out_to_MUX_Add123_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg725_out_to_MUX_Add123_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg943_out_to_MUX_Add123_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg804_out_to_MUX_Add123_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg803_out_to_MUX_Add123_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg803_out_to_MUX_Add123_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg606_out_to_MUX_Add123_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add123_1_impl_1_out);

   Delay1No149_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add123_1_impl_1_out,
                 Y => Delay1No149_out);

Delay1No150_out_to_Add123_2_impl_parent_implementedSystem_port_0_cast <= Delay1No150_out;
Delay1No151_out_to_Add123_2_impl_parent_implementedSystem_port_1_cast <= Delay1No151_out;
   Add123_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add123_2_impl_out,
                 X => Delay1No150_out_to_Add123_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No151_out_to_Add123_2_impl_parent_implementedSystem_port_1_cast);

SharedReg920_out_to_MUX_Add123_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg920_out;
SharedReg302_out_to_MUX_Add123_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg302_out;
SharedReg651_out_to_MUX_Add123_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg651_out;
SharedReg728_out_to_MUX_Add123_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg728_out;
SharedReg554_out_to_MUX_Add123_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg554_out;
SharedReg10_out_to_MUX_Add123_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg10_out;
SharedReg536_out_to_MUX_Add123_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg536_out;
Delay6No44_out_to_MUX_Add123_2_impl_0_parent_implementedSystem_port_8_cast <= Delay6No44_out;
SharedReg421_out_to_MUX_Add123_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg421_out;
SharedReg919_out_to_MUX_Add123_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg919_out;
SharedReg919_out_to_MUX_Add123_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg919_out;
SharedReg726_out_to_MUX_Add123_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg726_out;
   MUX_Add123_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg920_out_to_MUX_Add123_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg302_out_to_MUX_Add123_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg919_out_to_MUX_Add123_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg726_out_to_MUX_Add123_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg651_out_to_MUX_Add123_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg728_out_to_MUX_Add123_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg554_out_to_MUX_Add123_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg10_out_to_MUX_Add123_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg536_out_to_MUX_Add123_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay6No44_out_to_MUX_Add123_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg421_out_to_MUX_Add123_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg919_out_to_MUX_Add123_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add123_2_impl_0_out);

   Delay1No150_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add123_2_impl_0_out,
                 Y => Delay1No150_out);

SharedReg946_out_to_MUX_Add123_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg946_out;
SharedReg264_out_to_MUX_Add123_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg264_out;
SharedReg726_out_to_MUX_Add123_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg726_out;
SharedReg808_out_to_MUX_Add123_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg808_out;
SharedReg609_out_to_MUX_Add123_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg609_out;
SharedReg26_out_to_MUX_Add123_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg26_out;
SharedReg808_out_to_MUX_Add123_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg808_out;
SharedReg921_out_to_MUX_Add123_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg921_out;
SharedReg487_out_to_MUX_Add123_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg487_out;
SharedReg945_out_to_MUX_Add123_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg945_out;
SharedReg945_out_to_MUX_Add123_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg945_out;
SharedReg806_out_to_MUX_Add123_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg806_out;
   MUX_Add123_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg946_out_to_MUX_Add123_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg264_out_to_MUX_Add123_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg945_out_to_MUX_Add123_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg806_out_to_MUX_Add123_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg726_out_to_MUX_Add123_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg808_out_to_MUX_Add123_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg609_out_to_MUX_Add123_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg26_out_to_MUX_Add123_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg808_out_to_MUX_Add123_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg921_out_to_MUX_Add123_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg487_out_to_MUX_Add123_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg945_out_to_MUX_Add123_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add123_2_impl_1_out);

   Delay1No151_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add123_2_impl_1_out,
                 Y => Delay1No151_out);

Delay1No152_out_to_Add123_3_impl_parent_implementedSystem_port_0_cast <= Delay1No152_out;
Delay1No153_out_to_Add123_3_impl_parent_implementedSystem_port_1_cast <= Delay1No153_out;
   Add123_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add123_3_impl_out,
                 X => Delay1No152_out_to_Add123_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No153_out_to_Add123_3_impl_parent_implementedSystem_port_1_cast);

SharedReg730_out_to_MUX_Add123_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg730_out;
SharedReg923_out_to_MUX_Add123_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg923_out;
SharedReg266_out_to_MUX_Add123_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg266_out;
SharedReg192_out_to_MUX_Add123_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg192_out;
SharedReg732_out_to_MUX_Add123_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg732_out;
SharedReg556_out_to_MUX_Add123_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg556_out;
SharedReg6_out_to_MUX_Add123_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg6_out;
SharedReg539_out_to_MUX_Add123_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg539_out;
SharedReg924_out_to_MUX_Add123_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg924_out;
SharedReg423_out_to_MUX_Add123_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg423_out;
SharedReg923_out_to_MUX_Add123_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg923_out;
SharedReg923_out_to_MUX_Add123_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg923_out;
   MUX_Add123_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg730_out_to_MUX_Add123_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg923_out_to_MUX_Add123_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg923_out_to_MUX_Add123_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg923_out_to_MUX_Add123_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg266_out_to_MUX_Add123_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg192_out_to_MUX_Add123_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg732_out_to_MUX_Add123_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg556_out_to_MUX_Add123_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg6_out_to_MUX_Add123_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg539_out_to_MUX_Add123_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg924_out_to_MUX_Add123_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg423_out_to_MUX_Add123_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add123_3_impl_0_out);

   Delay1No152_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add123_3_impl_0_out,
                 Y => Delay1No152_out);

SharedReg809_out_to_MUX_Add123_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg809_out;
SharedReg948_out_to_MUX_Add123_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg948_out;
SharedReg247_out_to_MUX_Add123_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg247_out;
SharedReg353_out_to_MUX_Add123_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg353_out;
SharedReg811_out_to_MUX_Add123_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg811_out;
SharedReg612_out_to_MUX_Add123_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg612_out;
SharedReg22_out_to_MUX_Add123_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg22_out;
SharedReg811_out_to_MUX_Add123_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg811_out;
SharedReg949_out_to_MUX_Add123_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg949_out;
SharedReg490_out_to_MUX_Add123_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg490_out;
SharedReg948_out_to_MUX_Add123_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg948_out;
SharedReg948_out_to_MUX_Add123_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg948_out;
   MUX_Add123_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg809_out_to_MUX_Add123_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg948_out_to_MUX_Add123_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg948_out_to_MUX_Add123_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg948_out_to_MUX_Add123_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg247_out_to_MUX_Add123_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg353_out_to_MUX_Add123_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg811_out_to_MUX_Add123_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg612_out_to_MUX_Add123_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg22_out_to_MUX_Add123_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg811_out_to_MUX_Add123_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg949_out_to_MUX_Add123_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg490_out_to_MUX_Add123_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add123_3_impl_1_out);

   Delay1No153_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add123_3_impl_1_out,
                 Y => Delay1No153_out);

Delay1No154_out_to_Add123_6_impl_parent_implementedSystem_port_0_cast <= Delay1No154_out;
Delay1No155_out_to_Add123_6_impl_parent_implementedSystem_port_1_cast <= Delay1No155_out;
   Add123_6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add123_6_impl_out,
                 X => Delay1No154_out_to_Add123_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No155_out_to_Add123_6_impl_parent_implementedSystem_port_1_cast);

SharedReg847_out_to_MUX_Add123_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg847_out;
SharedReg936_out_to_MUX_Add123_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg936_out;
SharedReg429_out_to_MUX_Add123_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg429_out;
SharedReg742_out_to_MUX_Add123_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg742_out;
SharedReg742_out_to_MUX_Add123_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg742_out;
SharedReg562_out_to_MUX_Add123_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg562_out;
SharedReg525_out_to_MUX_Add123_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg525_out;
SharedReg320_out_to_MUX_Add123_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg320_out;
SharedReg382_out_to_MUX_Add123_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg382_out;
SharedReg935_out_to_MUX_Add123_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg935_out;
Delay4No223_out_to_MUX_Add123_6_impl_0_parent_implementedSystem_port_11_cast <= Delay4No223_out;
SharedReg10_out_to_MUX_Add123_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg10_out;
   MUX_Add123_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg847_out_to_MUX_Add123_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg936_out_to_MUX_Add123_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay4No223_out_to_MUX_Add123_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg10_out_to_MUX_Add123_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg429_out_to_MUX_Add123_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg742_out_to_MUX_Add123_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg742_out_to_MUX_Add123_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg562_out_to_MUX_Add123_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg525_out_to_MUX_Add123_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg320_out_to_MUX_Add123_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg382_out_to_MUX_Add123_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg935_out_to_MUX_Add123_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add123_6_impl_0_out);

   Delay1No154_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add123_6_impl_0_out,
                 Y => Delay1No154_out);

SharedReg643_out_to_MUX_Add123_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg643_out;
SharedReg958_out_to_MUX_Add123_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg958_out;
SharedReg499_out_to_MUX_Add123_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg499_out;
SharedReg818_out_to_MUX_Add123_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg818_out;
SharedReg818_out_to_MUX_Add123_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg818_out;
SharedReg621_out_to_MUX_Add123_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg621_out;
SharedReg547_out_to_MUX_Add123_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg547_out;
SharedReg324_out_to_MUX_Add123_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg324_out;
SharedReg387_out_to_MUX_Add123_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg387_out;
SharedReg908_out_to_MUX_Add123_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg908_out;
Delay4No230_out_to_MUX_Add123_6_impl_1_parent_implementedSystem_port_11_cast <= Delay4No230_out;
SharedReg26_out_to_MUX_Add123_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg26_out;
   MUX_Add123_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg643_out_to_MUX_Add123_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg958_out_to_MUX_Add123_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay4No230_out_to_MUX_Add123_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg26_out_to_MUX_Add123_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg499_out_to_MUX_Add123_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg818_out_to_MUX_Add123_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg818_out_to_MUX_Add123_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg621_out_to_MUX_Add123_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg547_out_to_MUX_Add123_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg324_out_to_MUX_Add123_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg387_out_to_MUX_Add123_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg908_out_to_MUX_Add123_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add123_6_impl_1_out);

   Delay1No155_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add123_6_impl_1_out,
                 Y => Delay1No155_out);

Delay1No156_out_to_Add35_0_impl_parent_implementedSystem_port_0_cast <= Delay1No156_out;
Delay1No157_out_to_Add35_0_impl_parent_implementedSystem_port_1_cast <= Delay1No157_out;
   Add35_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add35_0_impl_out,
                 X => Delay1No156_out_to_Add35_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No157_out_to_Add35_0_impl_parent_implementedSystem_port_1_cast);

SharedReg914_out_to_MUX_Add35_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg914_out;
SharedReg13_out_to_MUX_Add35_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg13_out;
SharedReg823_out_to_MUX_Add35_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg823_out;
Delay6No42_out_to_MUX_Add35_0_impl_0_parent_implementedSystem_port_4_cast <= Delay6No42_out;
SharedReg417_out_to_MUX_Add35_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg417_out;
SharedReg911_out_to_MUX_Add35_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg911_out;
SharedReg911_out_to_MUX_Add35_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg911_out;
SharedReg718_out_to_MUX_Add35_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg718_out;
SharedReg912_out_to_MUX_Add35_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg912_out;
SharedReg1037_out_to_MUX_Add35_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1037_out;
SharedReg626_out_to_MUX_Add35_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg626_out;
SharedReg961_out_to_MUX_Add35_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg961_out;
   MUX_Add35_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg914_out_to_MUX_Add35_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg13_out_to_MUX_Add35_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg626_out_to_MUX_Add35_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg961_out_to_MUX_Add35_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg823_out_to_MUX_Add35_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay6No42_out_to_MUX_Add35_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg417_out_to_MUX_Add35_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg911_out_to_MUX_Add35_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg911_out_to_MUX_Add35_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg718_out_to_MUX_Add35_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg912_out_to_MUX_Add35_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1037_out_to_MUX_Add35_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add35_0_impl_0_out);

   Delay1No156_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add35_0_impl_0_out,
                 Y => Delay1No156_out);

Delay4No259_out_to_MUX_Add35_0_impl_1_parent_implementedSystem_port_1_cast <= Delay4No259_out;
SharedReg29_out_to_MUX_Add35_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg29_out;
SharedReg625_out_to_MUX_Add35_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg625_out;
SharedReg913_out_to_MUX_Add35_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg913_out;
SharedReg481_out_to_MUX_Add35_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg481_out;
SharedReg939_out_to_MUX_Add35_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg939_out;
SharedReg939_out_to_MUX_Add35_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg939_out;
SharedReg800_out_to_MUX_Add35_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg800_out;
SharedReg940_out_to_MUX_Add35_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg940_out;
SharedReg1041_out_to_MUX_Add35_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1041_out;
SharedReg397_out_to_MUX_Add35_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg397_out;
SharedReg939_out_to_MUX_Add35_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg939_out;
   MUX_Add35_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay4No259_out_to_MUX_Add35_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg29_out_to_MUX_Add35_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg397_out_to_MUX_Add35_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg939_out_to_MUX_Add35_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg625_out_to_MUX_Add35_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg913_out_to_MUX_Add35_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg481_out_to_MUX_Add35_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg939_out_to_MUX_Add35_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg939_out_to_MUX_Add35_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg800_out_to_MUX_Add35_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg940_out_to_MUX_Add35_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1041_out_to_MUX_Add35_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add35_0_impl_1_out);

   Delay1No157_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add35_0_impl_1_out,
                 Y => Delay1No157_out);

Delay1No158_out_to_Add35_1_impl_parent_implementedSystem_port_0_cast <= Delay1No158_out;
Delay1No159_out_to_Add35_1_impl_parent_implementedSystem_port_1_cast <= Delay1No159_out;
   Add35_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add35_1_impl_out,
                 X => Delay1No158_out_to_Add35_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No159_out_to_Add35_1_impl_parent_implementedSystem_port_1_cast);

SharedReg629_out_to_MUX_Add35_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg629_out;
SharedReg915_out_to_MUX_Add35_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg915_out;
Delay4No218_out_to_MUX_Add35_1_impl_0_parent_implementedSystem_port_3_cast <= Delay4No218_out;
SharedReg10_out_to_MUX_Add35_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg10_out;
SharedReg533_out_to_MUX_Add35_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg533_out;
Delay6No43_out_to_MUX_Add35_1_impl_0_parent_implementedSystem_port_6_cast <= Delay6No43_out;
SharedReg419_out_to_MUX_Add35_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg419_out;
SharedReg915_out_to_MUX_Add35_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg915_out;
SharedReg915_out_to_MUX_Add35_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg915_out;
SharedReg722_out_to_MUX_Add35_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg722_out;
SharedReg916_out_to_MUX_Add35_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg916_out;
SharedReg1007_out_to_MUX_Add35_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1007_out;
   MUX_Add35_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg629_out_to_MUX_Add35_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg915_out_to_MUX_Add35_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg916_out_to_MUX_Add35_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1007_out_to_MUX_Add35_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => Delay4No218_out_to_MUX_Add35_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg10_out_to_MUX_Add35_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg533_out_to_MUX_Add35_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay6No43_out_to_MUX_Add35_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg419_out_to_MUX_Add35_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg915_out_to_MUX_Add35_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg915_out_to_MUX_Add35_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg722_out_to_MUX_Add35_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add35_1_impl_0_out);

   Delay1No158_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add35_1_impl_0_out,
                 Y => Delay1No158_out);

SharedReg400_out_to_MUX_Add35_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg400_out;
SharedReg888_out_to_MUX_Add35_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg888_out;
Delay4No225_out_to_MUX_Add35_1_impl_1_parent_implementedSystem_port_3_cast <= Delay4No225_out;
SharedReg26_out_to_MUX_Add35_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg26_out;
SharedReg805_out_to_MUX_Add35_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg805_out;
SharedReg917_out_to_MUX_Add35_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg917_out;
SharedReg484_out_to_MUX_Add35_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg484_out;
SharedReg942_out_to_MUX_Add35_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg942_out;
SharedReg942_out_to_MUX_Add35_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg942_out;
SharedReg803_out_to_MUX_Add35_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg803_out;
SharedReg943_out_to_MUX_Add35_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg943_out;
SharedReg1011_out_to_MUX_Add35_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1011_out;
   MUX_Add35_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg400_out_to_MUX_Add35_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg888_out_to_MUX_Add35_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg943_out_to_MUX_Add35_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1011_out_to_MUX_Add35_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => Delay4No225_out_to_MUX_Add35_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg26_out_to_MUX_Add35_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg805_out_to_MUX_Add35_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg917_out_to_MUX_Add35_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg484_out_to_MUX_Add35_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg942_out_to_MUX_Add35_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg942_out_to_MUX_Add35_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg803_out_to_MUX_Add35_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add35_1_impl_1_out);

   Delay1No159_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add35_1_impl_1_out,
                 Y => Delay1No159_out);

Delay1No160_out_to_Add35_6_impl_parent_implementedSystem_port_0_cast <= Delay1No160_out;
Delay1No161_out_to_Add35_6_impl_parent_implementedSystem_port_1_cast <= Delay1No161_out;
   Add35_6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add35_6_impl_out,
                 X => Delay1No160_out_to_Add35_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No161_out_to_Add35_6_impl_parent_implementedSystem_port_1_cast);

SharedReg743_out_to_MUX_Add35_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg743_out;
Delay6No48_out_to_MUX_Add35_6_impl_0_parent_implementedSystem_port_2_cast <= Delay6No48_out;
SharedReg936_out_to_MUX_Add35_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg936_out;
SharedReg935_out_to_MUX_Add35_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg935_out;
SharedReg935_out_to_MUX_Add35_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg935_out;
SharedReg742_out_to_MUX_Add35_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg742_out;
SharedReg935_out_to_MUX_Add35_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg935_out;
SharedReg1033_out_to_MUX_Add35_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1033_out;
SharedReg663_out_to_MUX_Add35_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg663_out;
SharedReg979_out_to_MUX_Add35_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg979_out;
SharedReg938_out_to_MUX_Add35_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg938_out;
SharedReg13_out_to_MUX_Add35_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg13_out;
   MUX_Add35_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg743_out_to_MUX_Add35_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay6No48_out_to_MUX_Add35_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg938_out_to_MUX_Add35_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg13_out_to_MUX_Add35_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg936_out_to_MUX_Add35_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg935_out_to_MUX_Add35_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg935_out_to_MUX_Add35_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg742_out_to_MUX_Add35_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg935_out_to_MUX_Add35_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1033_out_to_MUX_Add35_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg663_out_to_MUX_Add35_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg979_out_to_MUX_Add35_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add35_6_impl_0_out);

   Delay1No160_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add35_6_impl_0_out,
                 Y => Delay1No160_out);

SharedReg819_out_to_MUX_Add35_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg819_out;
SharedReg937_out_to_MUX_Add35_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg937_out;
SharedReg958_out_to_MUX_Add35_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg958_out;
SharedReg957_out_to_MUX_Add35_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg957_out;
SharedReg957_out_to_MUX_Add35_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg957_out;
SharedReg818_out_to_MUX_Add35_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg818_out;
SharedReg957_out_to_MUX_Add35_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg957_out;
SharedReg1069_out_to_MUX_Add35_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1069_out;
SharedReg742_out_to_MUX_Add35_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg742_out;
SharedReg957_out_to_MUX_Add35_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg957_out;
Delay4No265_out_to_MUX_Add35_6_impl_1_parent_implementedSystem_port_11_cast <= Delay4No265_out;
SharedReg29_out_to_MUX_Add35_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg29_out;
   MUX_Add35_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg819_out_to_MUX_Add35_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg937_out_to_MUX_Add35_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay4No265_out_to_MUX_Add35_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg29_out_to_MUX_Add35_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg958_out_to_MUX_Add35_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg957_out_to_MUX_Add35_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg957_out_to_MUX_Add35_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg818_out_to_MUX_Add35_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg957_out_to_MUX_Add35_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1069_out_to_MUX_Add35_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg742_out_to_MUX_Add35_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg957_out_to_MUX_Add35_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Add35_6_impl_1_out);

   Delay1No161_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add35_6_impl_1_out,
                 Y => Delay1No161_out);

Delay1No162_out_to_Add130_6_impl_parent_implementedSystem_port_0_cast <= Delay1No162_out;
Delay1No163_out_to_Add130_6_impl_parent_implementedSystem_port_1_cast <= Delay1No163_out;
   Add130_6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add130_6_impl_out,
                 X => Delay1No162_out_to_Add130_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No163_out_to_Add130_6_impl_parent_implementedSystem_port_1_cast);

SharedReg15_out_to_MUX_Add130_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg15_out;
SharedReg644_out_to_MUX_Add130_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg644_out;
SharedReg936_out_to_MUX_Add130_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg936_out;
SharedReg980_out_to_MUX_Add130_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg980_out;
   MUX_Add130_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg15_out_to_MUX_Add130_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg644_out_to_MUX_Add130_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg936_out_to_MUX_Add130_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg980_out_to_MUX_Add130_6_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => MUX_Add130_6_impl_0_LUT_out,
                 oMux => MUX_Add130_6_impl_0_out);

   Delay1No162_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add130_6_impl_0_out,
                 Y => Delay1No162_out);

SharedReg31_out_to_MUX_Add130_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg31_out;
SharedReg415_out_to_MUX_Add130_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg415_out;
SharedReg958_out_to_MUX_Add130_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg958_out;
SharedReg938_out_to_MUX_Add130_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg938_out;
   MUX_Add130_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg31_out_to_MUX_Add130_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg415_out_to_MUX_Add130_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg958_out_to_MUX_Add130_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg938_out_to_MUX_Add130_6_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => MUX_Add130_6_impl_1_LUT_out,
                 oMux => MUX_Add130_6_impl_1_out);

   Delay1No163_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add130_6_impl_1_out,
                 Y => Delay1No163_out);

Delay1No164_out_to_Product4_0_impl_parent_implementedSystem_port_0_cast <= Delay1No164_out;
Delay1No165_out_to_Product4_0_impl_parent_implementedSystem_port_1_cast <= Delay1No165_out;
   Product4_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_0_impl_out,
                 X => Delay1No164_out_to_Product4_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No165_out_to_Product4_0_impl_parent_implementedSystem_port_1_cast);

SharedReg1108_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1108_out;
SharedReg1109_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1109_out;
SharedReg1111_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1111_out;
SharedReg1112_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1112_out;
SharedReg1122_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1122_out;
SharedReg1114_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1114_out;
SharedReg1103_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1103_out;
SharedReg1104_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1104_out;
SharedReg982_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg982_out;
SharedReg1143_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1143_out;
SharedReg1107_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1113_out;
   MUX_Product4_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1108_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1109_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1107_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1113_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1111_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1112_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1122_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1114_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1103_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1104_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg982_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1143_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product4_0_impl_0_out);

   Delay1No164_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_0_impl_0_out,
                 Y => Delay1No164_out);

SharedReg202_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg202_out;
SharedReg249_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg249_out;
SharedReg65_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg65_out;
SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg32_out;
SharedReg68_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg68_out;
SharedReg37_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg37_out;
SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg32_out;
SharedReg66_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg66_out;
SharedReg1133_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1133_out;
SharedReg1072_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1072_out;
SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg32_out;
SharedReg67_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg67_out;
   MUX_Product4_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg202_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg249_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg67_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg65_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg68_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg37_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg66_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1133_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1072_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product4_0_impl_1_out);

   Delay1No165_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_0_impl_1_out,
                 Y => Delay1No165_out);

Delay1No166_out_to_Product4_1_impl_parent_implementedSystem_port_0_cast <= Delay1No166_out;
Delay1No167_out_to_Product4_1_impl_parent_implementedSystem_port_1_cast <= Delay1No167_out;
   Product4_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_1_impl_out,
                 X => Delay1No166_out_to_Product4_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No167_out_to_Product4_1_impl_parent_implementedSystem_port_1_cast);

SharedReg1107_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1113_out;
SharedReg1108_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1108_out;
SharedReg1109_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1109_out;
SharedReg1111_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1111_out;
SharedReg1112_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1112_out;
SharedReg1122_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1122_out;
SharedReg1114_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1114_out;
SharedReg1103_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1103_out;
SharedReg1104_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1104_out;
SharedReg985_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg985_out;
SharedReg1143_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1143_out;
   MUX_Product4_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1107_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1113_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg985_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1143_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1108_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1109_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1111_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1112_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1122_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1114_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1103_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1104_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product4_1_impl_0_out);

   Delay1No166_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_1_impl_0_out,
                 Y => Delay1No166_out);

SharedReg158_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg158_out;
SharedReg39_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg39_out;
SharedReg130_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg130_out;
SharedReg234_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg234_out;
SharedReg38_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg38_out;
SharedReg158_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg158_out;
SharedReg40_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg40_out;
SharedReg163_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg163_out;
SharedReg38_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg38_out;
SharedReg70_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg70_out;
SharedReg1133_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1133_out;
SharedReg1083_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1083_out;
   MUX_Product4_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg158_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg39_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1133_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1083_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg130_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg234_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg38_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg158_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg40_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg163_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg38_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg70_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product4_1_impl_1_out);

   Delay1No167_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_1_impl_1_out,
                 Y => Delay1No167_out);

Delay1No168_out_to_Product4_2_impl_parent_implementedSystem_port_0_cast <= Delay1No168_out;
Delay1No169_out_to_Product4_2_impl_parent_implementedSystem_port_1_cast <= Delay1No169_out;
   Product4_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_2_impl_out,
                 X => Delay1No168_out_to_Product4_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No169_out_to_Product4_2_impl_parent_implementedSystem_port_1_cast);

SharedReg859_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg859_out;
SharedReg1143_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1143_out;
SharedReg1107_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1113_out;
SharedReg1108_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1108_out;
SharedReg1109_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1109_out;
SharedReg1111_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1111_out;
SharedReg1112_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1112_out;
SharedReg1122_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1122_out;
SharedReg1114_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1114_out;
SharedReg1103_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1103_out;
SharedReg1104_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1104_out;
   MUX_Product4_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg859_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1143_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1103_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1104_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1107_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1113_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1108_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1109_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1111_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1112_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1122_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1114_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product4_2_impl_0_out);

   Delay1No168_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_2_impl_0_out,
                 Y => Delay1No168_out);

SharedReg1133_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1133_out;
SharedReg1049_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1049_out;
SharedReg164_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg164_out;
SharedReg42_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg42_out;
SharedReg134_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg134_out;
SharedReg239_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg239_out;
SharedReg73_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg73_out;
SharedReg41_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg41_out;
SharedReg43_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg43_out;
SharedReg169_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg169_out;
SharedReg41_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg41_out;
SharedReg74_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg74_out;
   MUX_Product4_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1133_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1049_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg41_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg74_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg164_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg42_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg134_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg239_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg73_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg41_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg43_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg169_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product4_2_impl_1_out);

   Delay1No169_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_2_impl_1_out,
                 Y => Delay1No169_out);

Delay1No170_out_to_Product4_3_impl_parent_implementedSystem_port_0_cast <= Delay1No170_out;
Delay1No171_out_to_Product4_3_impl_parent_implementedSystem_port_1_cast <= Delay1No171_out;
   Product4_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_3_impl_out,
                 X => Delay1No170_out_to_Product4_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No171_out_to_Product4_3_impl_parent_implementedSystem_port_1_cast);

SharedReg1104_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1104_out;
SharedReg862_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg862_out;
SharedReg1143_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1143_out;
SharedReg1107_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1113_out;
SharedReg1108_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1108_out;
SharedReg1109_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1109_out;
SharedReg1111_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1111_out;
SharedReg1112_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1112_out;
SharedReg1122_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1122_out;
SharedReg1114_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1114_out;
SharedReg1103_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1103_out;
   MUX_Product4_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1104_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg862_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1114_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1103_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1143_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1107_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1113_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1108_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1109_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1111_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1112_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1122_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product4_3_impl_0_out);

   Delay1No170_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_3_impl_0_out,
                 Y => Delay1No170_out);

SharedReg78_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg78_out;
SharedReg1133_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1133_out;
SharedReg1055_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1055_out;
SharedReg170_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg170_out;
SharedReg199_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg199_out;
SharedReg110_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg110_out;
SharedReg244_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg244_out;
SharedReg44_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg44_out;
SharedReg44_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg44_out;
SharedReg47_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg47_out;
SharedReg174_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg174_out;
SharedReg44_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg44_out;
   MUX_Product4_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg78_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1133_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg174_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg44_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1055_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg170_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg199_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg110_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg244_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg44_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg44_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg47_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product4_3_impl_1_out);

   Delay1No171_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_3_impl_1_out,
                 Y => Delay1No171_out);

Delay1No172_out_to_Product4_4_impl_parent_implementedSystem_port_0_cast <= Delay1No172_out;
Delay1No173_out_to_Product4_4_impl_parent_implementedSystem_port_1_cast <= Delay1No173_out;
   Product4_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_4_impl_out,
                 X => Delay1No172_out_to_Product4_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No173_out_to_Product4_4_impl_parent_implementedSystem_port_1_cast);

SharedReg1114_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1114_out;
SharedReg1103_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1103_out;
SharedReg1104_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1104_out;
SharedReg690_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg690_out;
SharedReg1143_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1143_out;
SharedReg1107_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1113_out;
SharedReg1108_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1108_out;
SharedReg1109_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1109_out;
SharedReg1111_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1111_out;
SharedReg1112_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1112_out;
SharedReg1122_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1122_out;
   MUX_Product4_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1114_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1103_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1112_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1122_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1104_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg690_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1143_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1107_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1113_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1108_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1109_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1111_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product4_4_impl_0_out);

   Delay1No172_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_4_impl_0_out,
                 Y => Delay1No172_out);

SharedReg196_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg196_out;
SharedReg48_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg48_out;
SharedReg82_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg82_out;
SharedReg1133_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1133_out;
SharedReg1023_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1023_out;
SharedReg191_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg191_out;
SharedReg177_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg177_out;
SharedReg145_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg145_out;
SharedReg272_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg272_out;
SharedReg81_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg81_out;
SharedReg48_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg48_out;
SharedReg84_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg84_out;
   MUX_Product4_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg196_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg48_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg48_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg84_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg82_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1133_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1023_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg191_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg177_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg145_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg272_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg81_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product4_4_impl_1_out);

   Delay1No173_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_4_impl_1_out,
                 Y => Delay1No173_out);

Delay1No174_out_to_Product4_5_impl_parent_implementedSystem_port_0_cast <= Delay1No174_out;
Delay1No175_out_to_Product4_5_impl_parent_implementedSystem_port_1_cast <= Delay1No175_out;
   Product4_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_5_impl_out,
                 X => Delay1No174_out_to_Product4_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No175_out_to_Product4_5_impl_parent_implementedSystem_port_1_cast);

SharedReg1112_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1112_out;
SharedReg1122_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1122_out;
SharedReg1114_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1114_out;
SharedReg1103_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1103_out;
SharedReg1104_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1104_out;
SharedReg695_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg695_out;
SharedReg1143_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1143_out;
SharedReg1107_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1113_out;
SharedReg1108_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1108_out;
SharedReg1109_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1109_out;
SharedReg1111_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1111_out;
   MUX_Product4_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1112_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1122_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1109_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1111_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1114_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1103_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1104_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg695_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1143_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1107_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1113_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1108_out_to_MUX_Product4_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product4_5_impl_0_out);

   Delay1No174_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_5_impl_0_out,
                 Y => Delay1No174_out);

SharedReg86_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg86_out;
SharedReg121_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg121_out;
SharedReg57_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg57_out;
SharedReg52_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg52_out;
SharedReg87_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg87_out;
SharedReg1133_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1133_out;
SharedReg1030_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1030_out;
SharedReg52_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg52_out;
SharedReg88_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg88_out;
SharedReg212_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg212_out;
SharedReg286_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg286_out;
SharedReg150_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg150_out;
   MUX_Product4_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg86_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg121_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg286_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg150_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg57_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg52_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg87_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1133_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1030_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg52_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg88_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg212_out_to_MUX_Product4_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product4_5_impl_1_out);

   Delay1No175_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_5_impl_1_out,
                 Y => Delay1No175_out);

Delay1No176_out_to_Product4_6_impl_parent_implementedSystem_port_0_cast <= Delay1No176_out;
Delay1No177_out_to_Product4_6_impl_parent_implementedSystem_port_1_cast <= Delay1No177_out;
   Product4_6_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_6_impl_out,
                 X => Delay1No176_out_to_Product4_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No177_out_to_Product4_6_impl_parent_implementedSystem_port_1_cast);

SharedReg1111_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1111_out;
SharedReg1112_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1112_out;
SharedReg1122_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1122_out;
SharedReg1114_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1114_out;
SharedReg1103_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1103_out;
SharedReg1104_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1104_out;
SharedReg872_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg872_out;
SharedReg1143_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1143_out;
SharedReg1107_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1113_out;
SharedReg1108_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1108_out;
SharedReg1109_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1109_out;
   MUX_Product4_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1111_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1112_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1108_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1109_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1122_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1114_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1103_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1104_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg872_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1143_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1107_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1113_out_to_MUX_Product4_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product4_6_impl_0_out);

   Delay1No176_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_6_impl_0_out,
                 Y => Delay1No176_out);

SharedReg91_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg91_out;
SharedReg91_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg91_out;
SharedReg125_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg125_out;
SharedReg229_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg229_out;
SharedReg60_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg60_out;
SharedReg92_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg92_out;
SharedReg1133_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1133_out;
SharedReg1068_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1068_out;
SharedReg60_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg60_out;
SharedReg62_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg62_out;
SharedReg187_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg187_out;
SharedReg320_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg320_out;
   MUX_Product4_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg91_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg91_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg187_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg320_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg125_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg229_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg60_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg92_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1133_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1068_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg60_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg62_out_to_MUX_Product4_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product4_6_impl_1_out);

   Delay1No177_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_6_impl_1_out,
                 Y => Delay1No177_out);

Delay1No178_out_to_Product21_0_impl_parent_implementedSystem_port_0_cast <= Delay1No178_out;
Delay1No179_out_to_Product21_0_impl_parent_implementedSystem_port_1_cast <= Delay1No179_out;
   Product21_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_0_impl_out,
                 X => Delay1No178_out_to_Product21_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No179_out_to_Product21_0_impl_parent_implementedSystem_port_1_cast);

SharedReg1108_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1108_out;
SharedReg1109_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1109_out;
SharedReg1111_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1111_out;
SharedReg1112_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1112_out;
SharedReg98_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg98_out;
SharedReg1114_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1114_out;
SharedReg1115_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1115_out;
SharedReg66_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg66_out;
SharedReg1132_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1132_out;
SharedReg1072_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1072_out;
SharedReg1107_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1113_out;
   MUX_Product21_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1108_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1109_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1107_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1113_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1111_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1112_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg98_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1114_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1115_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg66_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1132_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1072_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product21_0_impl_0_out);

   Delay1No178_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_0_impl_0_out,
                 Y => Delay1No178_out);

SharedReg249_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg249_out;
SharedReg128_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg128_out;
SharedReg95_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg95_out;
SharedReg65_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg65_out;
SharedReg1122_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1122_out;
SharedReg32_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg32_out;
SharedReg32_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg32_out;
SharedReg1116_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1116_out;
SharedReg1039_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1039_out;
SharedReg1145_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1145_out;
SharedReg65_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg65_out;
SharedReg98_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg98_out;
   MUX_Product21_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg249_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg128_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg65_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg98_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg95_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg65_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1122_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg32_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg32_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1116_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1039_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1145_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product21_0_impl_1_out);

   Delay1No179_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_0_impl_1_out,
                 Y => Delay1No179_out);

Delay1No180_out_to_Product21_1_impl_parent_implementedSystem_port_0_cast <= Delay1No180_out;
Delay1No181_out_to_Product21_1_impl_parent_implementedSystem_port_1_cast <= Delay1No181_out;
   Product21_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_1_impl_out,
                 X => Delay1No180_out_to_Product21_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No181_out_to_Product21_1_impl_parent_implementedSystem_port_1_cast);

SharedReg1107_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1113_out;
SharedReg1108_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1108_out;
SharedReg1109_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1109_out;
SharedReg1111_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1111_out;
SharedReg1112_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1112_out;
SharedReg72_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg72_out;
SharedReg1114_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1114_out;
SharedReg1115_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1115_out;
SharedReg70_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg70_out;
SharedReg1132_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1132_out;
SharedReg1083_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1083_out;
   MUX_Product21_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1107_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1113_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1132_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1083_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1108_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1109_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1111_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1112_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg72_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1114_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1115_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg70_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product21_1_impl_0_out);

   Delay1No180_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_1_impl_0_out,
                 Y => Delay1No180_out);

SharedReg38_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg38_out;
SharedReg72_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg72_out;
SharedReg234_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg234_out;
SharedReg101_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg101_out;
SharedReg69_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg69_out;
SharedReg38_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg38_out;
SharedReg1122_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1122_out;
SharedReg38_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg38_out;
SharedReg38_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg38_out;
SharedReg1116_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1116_out;
SharedReg1044_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1044_out;
SharedReg1145_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1145_out;
   MUX_Product21_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg38_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg72_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1044_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1145_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg234_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg101_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg69_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg38_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1122_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg38_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg38_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1116_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product21_1_impl_1_out);

   Delay1No181_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_1_impl_1_out,
                 Y => Delay1No181_out);

Delay1No182_out_to_Product21_2_impl_parent_implementedSystem_port_0_cast <= Delay1No182_out;
Delay1No183_out_to_Product21_2_impl_parent_implementedSystem_port_1_cast <= Delay1No183_out;
   Product21_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_2_impl_out,
                 X => Delay1No182_out_to_Product21_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No183_out_to_Product21_2_impl_parent_implementedSystem_port_1_cast);

SharedReg1132_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1132_out;
SharedReg1049_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1049_out;
SharedReg1107_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1113_out;
SharedReg1108_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1108_out;
SharedReg1109_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1109_out;
SharedReg1111_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1111_out;
SharedReg1112_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1112_out;
SharedReg76_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg76_out;
SharedReg1114_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1114_out;
SharedReg1115_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1115_out;
SharedReg74_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg74_out;
   MUX_Product21_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1132_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1049_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1115_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg74_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1107_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1113_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1108_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1109_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1111_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1112_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg76_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1114_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product21_2_impl_0_out);

   Delay1No182_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_2_impl_0_out,
                 Y => Delay1No182_out);

SharedReg1014_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1014_out;
SharedReg1145_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1145_out;
SharedReg41_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg41_out;
SharedReg76_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg76_out;
SharedReg239_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg239_out;
SharedReg106_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg106_out;
SharedReg105_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg105_out;
SharedReg73_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg73_out;
SharedReg1122_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1122_out;
SharedReg73_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg73_out;
SharedReg41_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg41_out;
SharedReg1116_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1116_out;
   MUX_Product21_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1014_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1145_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg41_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1116_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg41_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg76_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg239_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg106_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg105_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg73_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1122_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg73_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product21_2_impl_1_out);

   Delay1No183_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_2_impl_1_out,
                 Y => Delay1No183_out);

Delay1No184_out_to_Product21_3_impl_parent_implementedSystem_port_0_cast <= Delay1No184_out;
Delay1No185_out_to_Product21_3_impl_parent_implementedSystem_port_1_cast <= Delay1No185_out;
   Product21_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_3_impl_out,
                 X => Delay1No184_out_to_Product21_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No185_out_to_Product21_3_impl_parent_implementedSystem_port_1_cast);

SharedReg78_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg78_out;
SharedReg1132_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1132_out;
SharedReg1055_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1055_out;
SharedReg1107_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1113_out;
SharedReg1108_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1108_out;
SharedReg1109_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1109_out;
SharedReg1111_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1111_out;
SharedReg1112_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1112_out;
SharedReg80_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg80_out;
SharedReg1114_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1114_out;
SharedReg1115_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1115_out;
   MUX_Product21_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg78_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1132_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1114_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1115_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1055_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1107_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1113_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1108_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1109_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1111_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1112_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg80_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product21_3_impl_0_out);

   Delay1No184_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_3_impl_0_out,
                 Y => Delay1No184_out);

SharedReg1116_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1116_out;
SharedReg1055_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1055_out;
SharedReg1145_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1145_out;
SharedReg198_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg198_out;
SharedReg80_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg80_out;
SharedReg139_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg139_out;
SharedReg78_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg78_out;
SharedReg77_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg77_out;
SharedReg77_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg77_out;
SharedReg1122_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1122_out;
SharedReg44_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg44_out;
SharedReg44_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg44_out;
   MUX_Product21_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1116_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1055_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg44_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg44_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1145_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg198_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg80_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg139_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg78_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg77_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg77_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1122_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product21_3_impl_1_out);

   Delay1No185_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_3_impl_1_out,
                 Y => Delay1No185_out);

Delay1No186_out_to_Product21_4_impl_parent_implementedSystem_port_0_cast <= Delay1No186_out;
Delay1No187_out_to_Product21_4_impl_parent_implementedSystem_port_1_cast <= Delay1No187_out;
   Product21_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_4_impl_out,
                 X => Delay1No186_out_to_Product21_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No187_out_to_Product21_4_impl_parent_implementedSystem_port_1_cast);

SharedReg1114_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1114_out;
SharedReg1115_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1115_out;
SharedReg82_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg82_out;
SharedReg1132_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1132_out;
SharedReg1023_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1023_out;
SharedReg1107_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1113_out;
SharedReg1108_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1108_out;
SharedReg1109_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1109_out;
SharedReg1111_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1111_out;
SharedReg1112_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1112_out;
SharedReg116_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg116_out;
   MUX_Product21_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1114_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1115_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1112_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg116_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg82_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1132_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1023_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1107_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1113_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1108_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1109_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1111_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product21_4_impl_0_out);

   Delay1No186_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_4_impl_0_out,
                 Y => Delay1No186_out);

SharedReg48_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg48_out;
SharedReg48_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg48_out;
SharedReg1116_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1116_out;
SharedReg1023_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1023_out;
SharedReg1145_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1145_out;
SharedReg175_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg175_out;
SharedReg51_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg51_out;
SharedReg206_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg206_out;
SharedReg115_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg115_out;
SharedReg114_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg114_out;
SharedReg81_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg81_out;
SharedReg1122_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1122_out;
   MUX_Product21_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg48_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg48_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg81_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1122_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1116_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1023_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1145_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg175_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg51_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg206_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg115_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg114_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product21_4_impl_1_out);

   Delay1No187_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_4_impl_1_out,
                 Y => Delay1No187_out);

Delay1No188_out_to_Product21_5_impl_parent_implementedSystem_port_0_cast <= Delay1No188_out;
Delay1No189_out_to_Product21_5_impl_parent_implementedSystem_port_1_cast <= Delay1No189_out;
   Product21_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_5_impl_out,
                 X => Delay1No188_out_to_Product21_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No189_out_to_Product21_5_impl_parent_implementedSystem_port_1_cast);

SharedReg1112_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1112_out;
SharedReg152_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg152_out;
SharedReg1114_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1114_out;
SharedReg1115_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1115_out;
SharedReg87_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg87_out;
SharedReg1132_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1132_out;
SharedReg1030_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1030_out;
SharedReg1107_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1113_out;
SharedReg1108_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1108_out;
SharedReg1109_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1109_out;
SharedReg1111_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1111_out;
   MUX_Product21_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1112_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg152_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1109_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1111_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1114_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1115_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg87_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1132_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1030_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1107_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1113_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1108_out_to_MUX_Product21_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product21_5_impl_0_out);

   Delay1No188_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_5_impl_0_out,
                 Y => Delay1No188_out);

SharedReg118_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg118_out;
SharedReg1122_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1122_out;
SharedReg86_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg86_out;
SharedReg52_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg52_out;
SharedReg1116_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1116_out;
SharedReg999_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg999_out;
SharedReg1145_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1145_out;
SharedReg86_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg86_out;
SharedReg89_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg89_out;
SharedReg286_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg286_out;
SharedReg183_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg183_out;
SharedReg182_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg182_out;
   MUX_Product21_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg118_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1122_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg183_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg182_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg86_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg52_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1116_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg999_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1145_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg86_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg89_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg286_out_to_MUX_Product21_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product21_5_impl_1_out);

   Delay1No189_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_5_impl_1_out,
                 Y => Delay1No189_out);

Delay1No190_out_to_Product21_6_impl_parent_implementedSystem_port_0_cast <= Delay1No190_out;
Delay1No191_out_to_Product21_6_impl_parent_implementedSystem_port_1_cast <= Delay1No191_out;
   Product21_6_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_6_impl_out,
                 X => Delay1No190_out_to_Product21_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No191_out_to_Product21_6_impl_parent_implementedSystem_port_1_cast);

SharedReg1111_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1111_out;
SharedReg1112_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1112_out;
SharedReg156_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg156_out;
SharedReg1114_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1114_out;
SharedReg1115_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1115_out;
SharedReg92_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg92_out;
SharedReg1132_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1132_out;
SharedReg1068_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1068_out;
SharedReg1107_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1113_out;
SharedReg1108_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1108_out;
SharedReg1109_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1109_out;
   MUX_Product21_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1111_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1112_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1108_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1109_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg156_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1114_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1115_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg92_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1132_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1068_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1107_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1113_out_to_MUX_Product21_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product21_6_impl_0_out);

   Delay1No190_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_6_impl_0_out,
                 Y => Delay1No190_out);

SharedReg123_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg123_out;
SharedReg123_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg123_out;
SharedReg1122_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1122_out;
SharedReg60_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg60_out;
SharedReg60_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg60_out;
SharedReg1116_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1116_out;
SharedReg1068_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1068_out;
SharedReg1145_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1145_out;
SharedReg91_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg91_out;
SharedReg125_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg125_out;
SharedReg218_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg218_out;
SharedReg154_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg154_out;
   MUX_Product21_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg123_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg123_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg218_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg154_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1122_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg60_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg60_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1116_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1068_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1145_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg91_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg125_out_to_MUX_Product21_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product21_6_impl_1_out);

   Delay1No191_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_6_impl_1_out,
                 Y => Delay1No191_out);

Delay1No192_out_to_Subtract2_0_impl_parent_implementedSystem_port_0_cast <= Delay1No192_out;
Delay1No193_out_to_Subtract2_0_impl_parent_implementedSystem_port_1_cast <= Delay1No193_out;
   Subtract2_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_0_impl_out,
                 X => Delay1No192_out_to_Subtract2_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No193_out_to_Subtract2_0_impl_parent_implementedSystem_port_1_cast);

SharedReg416_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg416_out;
SharedReg_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg_out;
SharedReg647_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg647_out;
SharedReg482_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg482_out;
SharedReg395_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg395_out;
SharedReg395_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg395_out;
SharedReg395_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg395_out;
SharedReg395_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg395_out;
SharedReg480_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg480_out;
SharedReg604_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg604_out;
SharedReg624_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg624_out;
SharedReg396_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg396_out;
   MUX_Subtract2_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg416_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg624_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg396_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg647_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg482_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg395_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg395_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg395_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg395_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg480_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg604_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract2_0_impl_0_out);

   Delay1No192_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_0_impl_0_out,
                 Y => Delay1No192_out);

SharedReg395_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg395_out;
SharedReg16_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg16_out;
SharedReg417_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg417_out;
Delay6No7_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_4_cast <= Delay6No7_out;
SharedReg501_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg501_out;
SharedReg501_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg501_out;
SharedReg501_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg501_out;
SharedReg501_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg501_out;
SharedReg550_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg550_out;
SharedReg417_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg417_out;
SharedReg800_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg800_out;
SharedReg416_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg416_out;
   MUX_Subtract2_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg395_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg16_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg800_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg416_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg417_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay6No7_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg501_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg501_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg501_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg501_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg550_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg417_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract2_0_impl_1_out);

   Delay1No193_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_0_impl_1_out,
                 Y => Delay1No193_out);

Delay1No194_out_to_Subtract2_1_impl_parent_implementedSystem_port_0_cast <= Delay1No194_out;
Delay1No195_out_to_Subtract2_1_impl_parent_implementedSystem_port_1_cast <= Delay1No195_out;
   Subtract2_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_1_impl_out,
                 X => Delay1No194_out_to_Subtract2_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No195_out_to_Subtract2_1_impl_parent_implementedSystem_port_1_cast);

SharedReg776_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg776_out;
SharedReg399_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg399_out;
SharedReg418_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg418_out;
SharedReg_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg_out;
SharedReg650_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg650_out;
SharedReg399_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg399_out;
SharedReg532_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg532_out;
SharedReg532_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg532_out;
SharedReg532_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg532_out;
SharedReg532_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg532_out;
SharedReg887_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg887_out;
SharedReg438_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg438_out;
   MUX_Subtract2_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg776_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg399_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg887_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg438_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg418_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg650_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg399_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg532_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg532_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg532_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg532_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract2_1_impl_0_out);

   Delay1No194_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_1_impl_0_out,
                 Y => Delay1No194_out);

SharedReg438_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg438_out;
SharedReg418_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg418_out;
SharedReg398_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg398_out;
SharedReg16_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg16_out;
SharedReg419_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg419_out;
SharedReg506_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg506_out;
SharedReg627_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg627_out;
SharedReg627_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg627_out;
SharedReg627_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg627_out;
SharedReg627_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg627_out;
SharedReg963_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg963_out;
SharedReg571_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg571_out;
   MUX_Subtract2_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg438_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg418_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg963_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg571_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg398_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg16_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg419_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg506_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg627_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg627_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg627_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg627_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract2_1_impl_1_out);

   Delay1No195_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_1_impl_1_out,
                 Y => Delay1No195_out);

Delay1No196_out_to_Subtract2_2_impl_parent_implementedSystem_port_0_cast <= Delay1No196_out;
Delay1No197_out_to_Subtract2_2_impl_parent_implementedSystem_port_1_cast <= Delay1No197_out;
   Subtract2_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_2_impl_out,
                 X => Delay1No196_out_to_Subtract2_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No197_out_to_Subtract2_2_impl_parent_implementedSystem_port_1_cast);

SharedReg892_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg892_out;
SharedReg746_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg746_out;
SharedReg784_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg784_out;
SharedReg402_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg402_out;
SharedReg420_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg420_out;
SharedReg1_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1_out;
SharedReg728_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg728_out;
SharedReg536_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg536_out;
SharedReg651_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg651_out;
SharedReg651_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg651_out;
SharedReg1014_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1014_out;
SharedReg651_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg651_out;
   MUX_Subtract2_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg892_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg746_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1014_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg651_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg784_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg402_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg420_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg728_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg536_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg651_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg651_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract2_2_impl_0_out);

   Delay1No196_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_2_impl_0_out,
                 Y => Delay1No196_out);

SharedReg967_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg967_out;
SharedReg446_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg446_out;
SharedReg746_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg746_out;
SharedReg420_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg420_out;
SharedReg401_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg401_out;
SharedReg17_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg17_out;
SharedReg555_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg555_out;
SharedReg631_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg631_out;
SharedReg829_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg829_out;
SharedReg829_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg829_out;
SharedReg752_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg752_out;
SharedReg829_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg829_out;
   MUX_Subtract2_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg967_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg446_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg752_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg829_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg746_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg420_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg401_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg17_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg555_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg631_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg829_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg829_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract2_2_impl_1_out);

   Delay1No197_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_2_impl_1_out,
                 Y => Delay1No197_out);

Delay1No198_out_to_Subtract2_3_impl_parent_implementedSystem_port_0_cast <= Delay1No198_out;
Delay1No199_out_to_Subtract2_3_impl_parent_implementedSystem_port_1_cast <= Delay1No199_out;
   Subtract2_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_3_impl_out,
                 X => Delay1No198_out_to_Subtract2_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No199_out_to_Subtract2_3_impl_parent_implementedSystem_port_1_cast);

SharedReg654_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg654_out;
SharedReg895_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg895_out;
SharedReg753_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg753_out;
SharedReg633_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg633_out;
SharedReg405_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg405_out;
SharedReg422_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg422_out;
SharedReg_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg_out;
SharedReg732_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg732_out;
SharedReg405_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg405_out;
SharedReg654_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg654_out;
SharedReg654_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg654_out;
SharedReg1019_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1019_out;
   MUX_Subtract2_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg654_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg895_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg654_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1019_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg753_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg633_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg405_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg422_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg732_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg405_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg654_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract2_3_impl_0_out);

   Delay1No198_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_3_impl_0_out,
                 Y => Delay1No198_out);

SharedReg833_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg833_out;
SharedReg969_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg969_out;
SharedReg581_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg581_out;
SharedReg809_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg809_out;
SharedReg422_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg422_out;
SharedReg404_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg404_out;
SharedReg16_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg16_out;
SharedReg557_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg557_out;
SharedReg514_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg514_out;
SharedReg833_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg833_out;
SharedReg833_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg833_out;
SharedReg757_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg757_out;
   MUX_Subtract2_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg833_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg969_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg833_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg757_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg581_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg809_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg422_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg404_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg16_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg557_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg514_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg833_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract2_3_impl_1_out);

   Delay1No199_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_3_impl_1_out,
                 Y => Delay1No199_out);

Delay1No200_out_to_Subtract2_4_impl_parent_implementedSystem_port_0_cast <= Delay1No200_out;
Delay1No201_out_to_Subtract2_4_impl_parent_implementedSystem_port_1_cast <= Delay1No201_out;
   Subtract2_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_4_impl_out,
                 X => Delay1No200_out_to_Subtract2_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No201_out_to_Subtract2_4_impl_parent_implementedSystem_port_1_cast);

SharedReg899_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg899_out;
SharedReg1023_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1023_out;
SharedReg657_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg657_out;
SharedReg899_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg899_out;
SharedReg758_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg758_out;
SharedReg791_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg791_out;
SharedReg408_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg408_out;
SharedReg541_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg541_out;
SharedReg1_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1_out;
SharedReg658_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg658_out;
SharedReg658_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg658_out;
SharedReg899_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg899_out;
   MUX_Subtract2_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg899_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1023_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg658_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg899_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg657_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg899_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg758_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg791_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg408_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg541_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg658_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract2_4_impl_0_out);

   Delay1No200_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_4_impl_0_out,
                 Y => Delay1No200_out);

SharedReg972_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg972_out;
SharedReg711_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg711_out;
SharedReg837_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg837_out;
SharedReg972_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg972_out;
SharedReg706_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg706_out;
SharedReg758_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg758_out;
SharedReg424_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg424_out;
SharedReg636_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg636_out;
SharedReg17_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg17_out;
SharedReg838_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg838_out;
SharedReg838_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg838_out;
SharedReg972_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg972_out;
   MUX_Subtract2_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg972_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg711_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg838_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg972_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg837_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg972_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg706_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg758_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg424_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg636_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg17_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg838_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract2_4_impl_1_out);

   Delay1No201_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_4_impl_1_out,
                 Y => Delay1No201_out);

Delay1No202_out_to_Subtract2_5_impl_parent_implementedSystem_port_0_cast <= Delay1No202_out;
Delay1No203_out_to_Subtract2_5_impl_parent_implementedSystem_port_1_cast <= Delay1No203_out;
   Subtract2_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_5_impl_out,
                 X => Delay1No202_out_to_Subtract2_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No203_out_to_Subtract2_5_impl_parent_implementedSystem_port_1_cast);

SharedReg661_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg661_out;
SharedReg660_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg660_out;
SharedReg660_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg660_out;
SharedReg544_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg544_out;
SharedReg544_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg544_out;
SharedReg903_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg903_out;
SharedReg619_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg619_out;
SharedReg765_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg765_out;
SharedReg411_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg411_out;
SharedReg544_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg544_out;
SharedReg2_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg2_out;
SharedReg661_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg661_out;
   MUX_Subtract2_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg661_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg660_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg2_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg661_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg660_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg544_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg544_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg903_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg619_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg765_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg411_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg544_out_to_MUX_Subtract2_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract2_5_impl_0_out);

   Delay1No202_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_5_impl_0_out,
                 Y => Delay1No202_out);

SharedReg842_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg842_out;
SharedReg841_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg841_out;
SharedReg841_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg841_out;
SharedReg639_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg639_out;
SharedReg639_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg639_out;
SharedReg975_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg975_out;
SharedReg427_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg427_out;
SharedReg712_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg712_out;
SharedReg426_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg426_out;
SharedReg639_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg639_out;
SharedReg18_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg18_out;
SharedReg842_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg842_out;
   MUX_Subtract2_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg842_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg841_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg18_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg842_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg841_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg639_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg639_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg975_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg427_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg712_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg426_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg639_out_to_MUX_Subtract2_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract2_5_impl_1_out);

   Delay1No203_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_5_impl_1_out,
                 Y => Delay1No203_out);

Delay1No204_out_to_Subtract2_6_impl_parent_implementedSystem_port_0_cast <= Delay1No204_out;
Delay1No205_out_to_Subtract2_6_impl_parent_implementedSystem_port_1_cast <= Delay1No205_out;
   Subtract2_6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_6_impl_out,
                 X => Delay1No204_out_to_Subtract2_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No205_out_to_Subtract2_6_impl_parent_implementedSystem_port_1_cast);

SharedReg744_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg744_out;
SharedReg500_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg500_out;
SharedReg547_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg547_out;
SharedReg413_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg413_out;
SharedReg413_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg413_out;
SharedReg413_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg413_out;
SharedReg290_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg290_out;
SharedReg622_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg622_out;
SharedReg217_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg217_out;
SharedReg414_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg414_out;
SharedReg428_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg428_out;
SharedReg_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg_out;
   MUX_Subtract2_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg744_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg500_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg428_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg547_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg413_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg413_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg413_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg290_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg622_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg217_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg414_out_to_MUX_Subtract2_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract2_6_impl_0_out);

   Delay1No204_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_6_impl_0_out,
                 Y => Delay1No204_out);

SharedReg563_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg563_out;
Delay6No13_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_2_cast <= Delay6No13_out;
SharedReg642_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg642_out;
SharedReg525_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg525_out;
SharedReg525_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg525_out;
SharedReg525_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg525_out;
SharedReg295_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg295_out;
SharedReg429_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg429_out;
SharedReg229_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg229_out;
SharedReg428_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg428_out;
SharedReg413_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg413_out;
SharedReg16_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg16_out;
   MUX_Subtract2_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg563_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay6No13_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg413_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg16_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg642_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg525_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg525_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg525_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg295_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg429_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg229_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg428_out_to_MUX_Subtract2_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract2_6_impl_1_out);

   Delay1No205_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_6_impl_1_out,
                 Y => Delay1No205_out);

Delay1No206_out_to_Product5_0_impl_parent_implementedSystem_port_0_cast <= Delay1No206_out;
Delay1No207_out_to_Product5_0_impl_parent_implementedSystem_port_1_cast <= Delay1No207_out;
   Product5_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product5_0_impl_out,
                 X => Delay1No206_out_to_Product5_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No207_out_to_Product5_0_impl_parent_implementedSystem_port_1_cast);

SharedReg1120_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1120_out;
SharedReg1121_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1121_out;
SharedReg1123_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1123_out;
SharedReg1124_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1124_out;
SharedReg1110_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1110_out;
SharedReg1126_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1126_out;
SharedReg1127_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1127_out;
SharedReg1104_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1104_out;
SharedReg1132_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1132_out;
SharedReg1147_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1147_out;
SharedReg1119_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1125_out;
   MUX_Product5_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1120_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1121_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1119_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1125_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1123_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1124_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1110_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1126_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1127_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1104_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1132_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1147_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product5_0_impl_0_out);

   Delay1No206_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product5_0_impl_0_out,
                 Y => Delay1No206_out);

SharedReg202_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg202_out;
SharedReg249_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg249_out;
SharedReg65_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg65_out;
SharedReg32_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg32_out;
SharedReg204_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg204_out;
SharedReg37_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg37_out;
SharedReg1004_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1004_out;
SharedReg96_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg96_out;
SharedReg982_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg982_out;
SharedReg1096_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1096_out;
SharedReg32_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg32_out;
SharedReg67_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg67_out;
   MUX_Product5_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg202_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg249_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg32_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg67_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg65_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg32_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg204_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg37_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1004_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg96_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg982_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1096_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product5_0_impl_1_out);

   Delay1No207_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product5_0_impl_1_out,
                 Y => Delay1No207_out);

Delay1No208_out_to_Product5_1_impl_parent_implementedSystem_port_0_cast <= Delay1No208_out;
Delay1No209_out_to_Product5_1_impl_parent_implementedSystem_port_1_cast <= Delay1No209_out;
   Product5_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product5_1_impl_out,
                 X => Delay1No208_out_to_Product5_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No209_out_to_Product5_1_impl_parent_implementedSystem_port_1_cast);

SharedReg1119_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1125_out;
SharedReg1120_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1120_out;
SharedReg1121_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1121_out;
SharedReg1123_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1123_out;
SharedReg1124_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1124_out;
SharedReg1110_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1110_out;
SharedReg1126_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1126_out;
SharedReg1127_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1127_out;
SharedReg1104_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1104_out;
SharedReg1132_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1132_out;
SharedReg1147_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1147_out;
   MUX_Product5_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1119_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1125_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1132_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1147_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1120_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1121_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1123_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1124_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1110_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1126_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1127_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1104_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product5_1_impl_0_out);

   Delay1No208_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product5_1_impl_0_out,
                 Y => Delay1No208_out);

SharedReg158_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg158_out;
SharedReg39_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg39_out;
SharedReg130_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg130_out;
SharedReg234_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg234_out;
SharedReg38_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg38_out;
SharedReg158_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg158_out;
SharedReg132_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg132_out;
SharedReg163_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg163_out;
SharedReg1007_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1007_out;
SharedReg101_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg101_out;
SharedReg985_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg985_out;
SharedReg785_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg785_out;
   MUX_Product5_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg158_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg39_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg985_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg785_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg130_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg234_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg38_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg158_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg132_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg163_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1007_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg101_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product5_1_impl_1_out);

   Delay1No209_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product5_1_impl_1_out,
                 Y => Delay1No209_out);

Delay1No210_out_to_Product5_2_impl_parent_implementedSystem_port_0_cast <= Delay1No210_out;
Delay1No211_out_to_Product5_2_impl_parent_implementedSystem_port_1_cast <= Delay1No211_out;
   Product5_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product5_2_impl_out,
                 X => Delay1No210_out_to_Product5_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No211_out_to_Product5_2_impl_parent_implementedSystem_port_1_cast);

SharedReg1132_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1132_out;
SharedReg1147_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1147_out;
SharedReg1119_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1125_out;
SharedReg1120_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1120_out;
SharedReg1121_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1121_out;
SharedReg1123_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1123_out;
SharedReg1124_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1124_out;
SharedReg1110_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1110_out;
SharedReg1126_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1126_out;
SharedReg1127_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1127_out;
SharedReg1104_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1104_out;
   MUX_Product5_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1132_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1147_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1127_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1104_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1119_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1125_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1120_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1121_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1123_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1124_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1110_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1126_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product5_2_impl_0_out);

   Delay1No210_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product5_2_impl_0_out,
                 Y => Delay1No210_out);

SharedReg859_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg859_out;
SharedReg878_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg878_out;
SharedReg164_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg164_out;
SharedReg42_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg42_out;
SharedReg134_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg134_out;
SharedReg239_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg239_out;
SharedReg73_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg73_out;
SharedReg41_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg41_out;
SharedReg136_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg136_out;
SharedReg169_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg169_out;
SharedReg986_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg986_out;
SharedReg106_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg106_out;
   MUX_Product5_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg859_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg878_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg986_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg106_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg164_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg42_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg134_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg239_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg73_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg41_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg136_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg169_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product5_2_impl_1_out);

   Delay1No211_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product5_2_impl_1_out,
                 Y => Delay1No211_out);

Delay1No212_out_to_Product5_3_impl_parent_implementedSystem_port_0_cast <= Delay1No212_out;
Delay1No213_out_to_Product5_3_impl_parent_implementedSystem_port_1_cast <= Delay1No213_out;
   Product5_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product5_3_impl_out,
                 X => Delay1No212_out_to_Product5_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No213_out_to_Product5_3_impl_parent_implementedSystem_port_1_cast);

SharedReg1104_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1104_out;
SharedReg1132_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1132_out;
SharedReg1147_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1147_out;
SharedReg1119_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1125_out;
SharedReg1120_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1120_out;
SharedReg1121_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1121_out;
SharedReg1123_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1123_out;
SharedReg1124_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1124_out;
SharedReg1110_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1110_out;
SharedReg1126_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1126_out;
SharedReg1127_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1127_out;
   MUX_Product5_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1104_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1132_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1126_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1127_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1147_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1119_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1125_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1120_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1121_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1123_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1124_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1110_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product5_3_impl_0_out);

   Delay1No212_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product5_3_impl_0_out,
                 Y => Delay1No212_out);

SharedReg111_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg111_out;
SharedReg862_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg862_out;
SharedReg792_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg792_out;
SharedReg170_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg170_out;
SharedReg199_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg199_out;
SharedReg110_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg110_out;
SharedReg244_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg244_out;
SharedReg44_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg44_out;
SharedReg44_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg44_out;
SharedReg142_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg142_out;
SharedReg174_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg174_out;
SharedReg1017_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1017_out;
   MUX_Product5_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg111_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg862_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg174_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1017_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg792_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg170_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg199_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg110_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg244_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg44_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg44_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg142_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product5_3_impl_1_out);

   Delay1No213_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product5_3_impl_1_out,
                 Y => Delay1No213_out);

Delay1No214_out_to_Product5_4_impl_parent_implementedSystem_port_0_cast <= Delay1No214_out;
Delay1No215_out_to_Product5_4_impl_parent_implementedSystem_port_1_cast <= Delay1No215_out;
   Product5_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product5_4_impl_out,
                 X => Delay1No214_out_to_Product5_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No215_out_to_Product5_4_impl_parent_implementedSystem_port_1_cast);

SharedReg1126_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1126_out;
SharedReg1127_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1127_out;
SharedReg1104_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1104_out;
SharedReg1132_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1132_out;
SharedReg1147_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1147_out;
SharedReg1119_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1125_out;
SharedReg1120_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1120_out;
SharedReg1121_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1121_out;
SharedReg1123_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1123_out;
SharedReg1124_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1124_out;
SharedReg1110_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1110_out;
   MUX_Product5_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1126_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1127_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1124_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1110_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1104_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1132_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1147_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1119_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1125_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1120_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1121_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1123_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product5_4_impl_0_out);

   Delay1No214_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product5_4_impl_0_out,
                 Y => Delay1No214_out);

SharedReg196_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg196_out;
SharedReg993_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg993_out;
SharedReg115_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg115_out;
SharedReg690_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg690_out;
SharedReg797_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg797_out;
SharedReg191_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg191_out;
SharedReg177_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg177_out;
SharedReg145_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg145_out;
SharedReg272_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg272_out;
SharedReg81_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg81_out;
SharedReg48_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg48_out;
SharedReg209_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg209_out;
   MUX_Product5_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg196_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg993_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg48_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg209_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg115_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg690_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg797_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg191_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg177_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg145_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg272_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg81_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product5_4_impl_1_out);

   Delay1No215_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product5_4_impl_1_out,
                 Y => Delay1No215_out);

Delay1No216_out_to_Product5_5_impl_parent_implementedSystem_port_0_cast <= Delay1No216_out;
Delay1No217_out_to_Product5_5_impl_parent_implementedSystem_port_1_cast <= Delay1No217_out;
   Product5_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product5_5_impl_out,
                 X => Delay1No216_out_to_Product5_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No217_out_to_Product5_5_impl_parent_implementedSystem_port_1_cast);

SharedReg1124_out_to_MUX_Product5_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1124_out;
SharedReg1110_out_to_MUX_Product5_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1110_out;
SharedReg1126_out_to_MUX_Product5_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1126_out;
SharedReg1127_out_to_MUX_Product5_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1127_out;
SharedReg1104_out_to_MUX_Product5_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1104_out;
SharedReg1132_out_to_MUX_Product5_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1132_out;
SharedReg1147_out_to_MUX_Product5_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1147_out;
SharedReg1119_out_to_MUX_Product5_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product5_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1125_out;
SharedReg1120_out_to_MUX_Product5_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1120_out;
SharedReg1121_out_to_MUX_Product5_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1121_out;
SharedReg1123_out_to_MUX_Product5_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1123_out;
   MUX_Product5_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1124_out_to_MUX_Product5_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1110_out_to_MUX_Product5_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1121_out_to_MUX_Product5_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1123_out_to_MUX_Product5_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1126_out_to_MUX_Product5_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1127_out_to_MUX_Product5_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1104_out_to_MUX_Product5_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1132_out_to_MUX_Product5_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1147_out_to_MUX_Product5_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1119_out_to_MUX_Product5_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1125_out_to_MUX_Product5_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1120_out_to_MUX_Product5_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product5_5_impl_0_out);

   Delay1No216_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product5_5_impl_0_out,
                 Y => Delay1No216_out);

SharedReg86_out_to_MUX_Product5_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg86_out;
SharedReg215_out_to_MUX_Product5_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg215_out;
SharedReg57_out_to_MUX_Product5_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg57_out;
SharedReg868_out_to_MUX_Product5_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg868_out;
SharedReg119_out_to_MUX_Product5_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg119_out;
SharedReg695_out_to_MUX_Product5_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg695_out;
SharedReg1061_out_to_MUX_Product5_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1061_out;
SharedReg52_out_to_MUX_Product5_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg52_out;
SharedReg88_out_to_MUX_Product5_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg88_out;
SharedReg212_out_to_MUX_Product5_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg212_out;
SharedReg286_out_to_MUX_Product5_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg286_out;
SharedReg150_out_to_MUX_Product5_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg150_out;
   MUX_Product5_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg86_out_to_MUX_Product5_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg215_out_to_MUX_Product5_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg286_out_to_MUX_Product5_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg150_out_to_MUX_Product5_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg57_out_to_MUX_Product5_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg868_out_to_MUX_Product5_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg119_out_to_MUX_Product5_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg695_out_to_MUX_Product5_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1061_out_to_MUX_Product5_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg52_out_to_MUX_Product5_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg88_out_to_MUX_Product5_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg212_out_to_MUX_Product5_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product5_5_impl_1_out);

   Delay1No217_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product5_5_impl_1_out,
                 Y => Delay1No217_out);

Delay1No218_out_to_Product5_6_impl_parent_implementedSystem_port_0_cast <= Delay1No218_out;
Delay1No219_out_to_Product5_6_impl_parent_implementedSystem_port_1_cast <= Delay1No219_out;
   Product5_6_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product5_6_impl_out,
                 X => Delay1No218_out_to_Product5_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No219_out_to_Product5_6_impl_parent_implementedSystem_port_1_cast);

SharedReg1123_out_to_MUX_Product5_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1123_out;
SharedReg1124_out_to_MUX_Product5_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1124_out;
SharedReg1110_out_to_MUX_Product5_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1110_out;
SharedReg1126_out_to_MUX_Product5_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1126_out;
SharedReg1127_out_to_MUX_Product5_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1127_out;
SharedReg1104_out_to_MUX_Product5_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1104_out;
SharedReg1132_out_to_MUX_Product5_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1132_out;
SharedReg1147_out_to_MUX_Product5_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1147_out;
SharedReg1119_out_to_MUX_Product5_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product5_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1125_out;
SharedReg1120_out_to_MUX_Product5_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1120_out;
SharedReg1121_out_to_MUX_Product5_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1121_out;
   MUX_Product5_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1123_out_to_MUX_Product5_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1124_out_to_MUX_Product5_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1120_out_to_MUX_Product5_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1121_out_to_MUX_Product5_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1110_out_to_MUX_Product5_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1126_out_to_MUX_Product5_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1127_out_to_MUX_Product5_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1104_out_to_MUX_Product5_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1132_out_to_MUX_Product5_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1147_out_to_MUX_Product5_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1119_out_to_MUX_Product5_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1125_out_to_MUX_Product5_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product5_6_impl_0_out);

   Delay1No218_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product5_6_impl_0_out,
                 Y => Delay1No218_out);

SharedReg91_out_to_MUX_Product5_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg91_out;
SharedReg91_out_to_MUX_Product5_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg91_out;
SharedReg221_out_to_MUX_Product5_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg221_out;
SharedReg229_out_to_MUX_Product5_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg229_out;
SharedReg1033_out_to_MUX_Product5_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1033_out;
SharedReg124_out_to_MUX_Product5_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg124_out;
SharedReg872_out_to_MUX_Product5_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg872_out;
SharedReg1077_out_to_MUX_Product5_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1077_out;
SharedReg60_out_to_MUX_Product5_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg60_out;
SharedReg62_out_to_MUX_Product5_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg62_out;
SharedReg187_out_to_MUX_Product5_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg187_out;
SharedReg320_out_to_MUX_Product5_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg320_out;
   MUX_Product5_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg91_out_to_MUX_Product5_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg91_out_to_MUX_Product5_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg187_out_to_MUX_Product5_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg320_out_to_MUX_Product5_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg221_out_to_MUX_Product5_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg229_out_to_MUX_Product5_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1033_out_to_MUX_Product5_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg124_out_to_MUX_Product5_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg872_out_to_MUX_Product5_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1077_out_to_MUX_Product5_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg60_out_to_MUX_Product5_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg62_out_to_MUX_Product5_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product5_6_impl_1_out);

   Delay1No219_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product5_6_impl_1_out,
                 Y => Delay1No219_out);

Delay1No220_out_to_Product12_0_impl_parent_implementedSystem_port_0_cast <= Delay1No220_out;
Delay1No221_out_to_Product12_0_impl_parent_implementedSystem_port_1_cast <= Delay1No221_out;
   Product12_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product12_0_impl_out,
                 X => Delay1No220_out_to_Product12_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No221_out_to_Product12_0_impl_parent_implementedSystem_port_1_cast);

SharedReg249_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg249_out;
SharedReg128_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg128_out;
SharedReg95_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg95_out;
SharedReg65_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg65_out;
SharedReg1110_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1110_out;
SharedReg32_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg32_out;
SharedReg1146_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1146_out;
SharedReg1104_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1104_out;
SharedReg1133_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1133_out;
SharedReg1151_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1151_out;
SharedReg65_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg65_out;
SharedReg98_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg98_out;
   MUX_Product12_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg249_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg128_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg65_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg98_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg95_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg65_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1110_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg32_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1146_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1104_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1133_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1151_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product12_0_impl_0_out);

   Delay1No220_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_0_impl_0_out,
                 Y => Delay1No220_out);

SharedReg1120_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1120_out;
SharedReg1121_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1121_out;
SharedReg1123_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1123_out;
SharedReg1124_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1124_out;
SharedReg35_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg35_out;
SharedReg1126_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1126_out;
SharedReg1094_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1094_out;
SharedReg128_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg128_out;
SharedReg1039_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1039_out;
SharedReg1096_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1096_out;
SharedReg1119_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1125_out;
   MUX_Product12_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1120_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1121_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1119_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1125_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1123_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1124_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg35_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1126_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1094_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg128_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1039_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1096_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product12_0_impl_1_out);

   Delay1No221_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_0_impl_1_out,
                 Y => Delay1No221_out);

Delay1No222_out_to_Product12_1_impl_parent_implementedSystem_port_0_cast <= Delay1No222_out;
Delay1No223_out_to_Product12_1_impl_parent_implementedSystem_port_1_cast <= Delay1No223_out;
   Product12_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product12_1_impl_out,
                 X => Delay1No222_out_to_Product12_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No223_out_to_Product12_1_impl_parent_implementedSystem_port_1_cast);

SharedReg38_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg38_out;
SharedReg72_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg72_out;
SharedReg234_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg234_out;
SharedReg101_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg101_out;
SharedReg69_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg69_out;
SharedReg38_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg38_out;
SharedReg1110_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1110_out;
SharedReg38_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg38_out;
SharedReg1146_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1146_out;
SharedReg1104_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1104_out;
SharedReg1133_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1133_out;
SharedReg1151_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1151_out;
   MUX_Product12_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg38_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg72_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1133_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1151_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg234_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg101_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg69_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg38_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1110_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg38_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1146_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1104_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product12_1_impl_0_out);

   Delay1No222_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_1_impl_0_out,
                 Y => Delay1No222_out);

SharedReg1119_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1125_out;
SharedReg1120_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1120_out;
SharedReg1121_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1121_out;
SharedReg1123_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1123_out;
SharedReg1124_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1124_out;
SharedReg161_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg161_out;
SharedReg1126_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1126_out;
SharedReg783_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg783_out;
SharedReg131_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg131_out;
SharedReg1044_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1044_out;
SharedReg785_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg785_out;
   MUX_Product12_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1119_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1125_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1044_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg785_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1120_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1121_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1123_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1124_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg161_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1126_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg783_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg131_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product12_1_impl_1_out);

   Delay1No223_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_1_impl_1_out,
                 Y => Delay1No223_out);

Delay1No224_out_to_Product12_2_impl_parent_implementedSystem_port_0_cast <= Delay1No224_out;
Delay1No225_out_to_Product12_2_impl_parent_implementedSystem_port_1_cast <= Delay1No225_out;
   Product12_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product12_2_impl_out,
                 X => Delay1No224_out_to_Product12_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No225_out_to_Product12_2_impl_parent_implementedSystem_port_1_cast);

SharedReg1133_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1133_out;
SharedReg1151_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1151_out;
SharedReg41_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg41_out;
SharedReg76_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg76_out;
SharedReg239_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg239_out;
SharedReg106_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg106_out;
SharedReg105_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg105_out;
SharedReg73_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg73_out;
SharedReg1110_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1110_out;
SharedReg73_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg73_out;
SharedReg1146_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1146_out;
SharedReg1104_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1104_out;
   MUX_Product12_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1133_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1151_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1146_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1104_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg41_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg76_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg239_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg106_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg105_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg73_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1110_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg73_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product12_2_impl_0_out);

   Delay1No224_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_2_impl_0_out,
                 Y => Delay1No224_out);

SharedReg1014_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1014_out;
SharedReg878_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg878_out;
SharedReg1119_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1125_out;
SharedReg1120_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1120_out;
SharedReg1121_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1121_out;
SharedReg1123_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1123_out;
SharedReg1124_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1124_out;
SharedReg166_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg166_out;
SharedReg1126_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1126_out;
SharedReg876_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg876_out;
SharedReg135_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg135_out;
   MUX_Product12_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1014_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg878_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg876_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg135_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1119_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1125_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1120_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1121_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1123_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1124_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg166_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1126_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product12_2_impl_1_out);

   Delay1No225_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_2_impl_1_out,
                 Y => Delay1No225_out);

Delay1No226_out_to_Product12_3_impl_parent_implementedSystem_port_0_cast <= Delay1No226_out;
Delay1No227_out_to_Product12_3_impl_parent_implementedSystem_port_1_cast <= Delay1No227_out;
   Product12_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product12_3_impl_out,
                 X => Delay1No226_out_to_Product12_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No227_out_to_Product12_3_impl_parent_implementedSystem_port_1_cast);

SharedReg1104_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1104_out;
SharedReg1133_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1133_out;
SharedReg1151_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1151_out;
SharedReg198_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg198_out;
SharedReg80_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg80_out;
SharedReg139_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg139_out;
SharedReg78_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg78_out;
SharedReg77_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg77_out;
SharedReg77_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg77_out;
SharedReg1110_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1110_out;
SharedReg44_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg44_out;
SharedReg1146_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1146_out;
   MUX_Product12_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1104_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1133_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg44_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1146_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1151_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg198_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg80_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg139_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg78_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg77_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg77_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1110_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product12_3_impl_0_out);

   Delay1No226_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_3_impl_0_out,
                 Y => Delay1No226_out);

SharedReg140_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg140_out;
SharedReg1055_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1055_out;
SharedReg792_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg792_out;
SharedReg1119_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1125_out;
SharedReg1120_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1120_out;
SharedReg1121_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1121_out;
SharedReg1123_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1123_out;
SharedReg1124_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1124_out;
SharedReg200_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg200_out;
SharedReg1126_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1126_out;
SharedReg758_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg758_out;
   MUX_Product12_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg140_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1055_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1126_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg758_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg792_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1119_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1125_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1120_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1121_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1123_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1124_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg200_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product12_3_impl_1_out);

   Delay1No227_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_3_impl_1_out,
                 Y => Delay1No227_out);

Delay1No228_out_to_Product12_4_impl_parent_implementedSystem_port_0_cast <= Delay1No228_out;
Delay1No229_out_to_Product12_4_impl_parent_implementedSystem_port_1_cast <= Delay1No229_out;
   Product12_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product12_4_impl_out,
                 X => Delay1No228_out_to_Product12_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No229_out_to_Product12_4_impl_parent_implementedSystem_port_1_cast);

SharedReg48_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg48_out;
SharedReg1146_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1146_out;
SharedReg1104_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1104_out;
SharedReg1133_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1133_out;
SharedReg1151_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1151_out;
SharedReg175_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg175_out;
SharedReg51_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg51_out;
SharedReg206_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg206_out;
SharedReg115_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg115_out;
SharedReg114_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg114_out;
SharedReg81_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg81_out;
SharedReg1110_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1110_out;
   MUX_Product12_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg48_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1146_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg81_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1110_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1104_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1133_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1151_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg175_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg51_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg206_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg115_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg114_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product12_4_impl_0_out);

   Delay1No228_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_4_impl_0_out,
                 Y => Delay1No228_out);

SharedReg1126_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1126_out;
SharedReg764_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg764_out;
SharedReg146_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg146_out;
SharedReg1023_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1023_out;
SharedReg797_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg797_out;
SharedReg1119_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1125_out;
SharedReg1120_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1120_out;
SharedReg1121_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1121_out;
SharedReg1123_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1123_out;
SharedReg1124_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1124_out;
SharedReg51_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg51_out;
   MUX_Product12_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1126_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg764_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1124_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg51_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg146_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1023_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg797_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1119_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1125_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1120_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1121_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1123_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product12_4_impl_1_out);

   Delay1No229_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_4_impl_1_out,
                 Y => Delay1No229_out);

Delay1No230_out_to_Product12_5_impl_parent_implementedSystem_port_0_cast <= Delay1No230_out;
Delay1No231_out_to_Product12_5_impl_parent_implementedSystem_port_1_cast <= Delay1No231_out;
   Product12_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product12_5_impl_out,
                 X => Delay1No230_out_to_Product12_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No231_out_to_Product12_5_impl_parent_implementedSystem_port_1_cast);

SharedReg118_out_to_MUX_Product12_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg118_out;
SharedReg1110_out_to_MUX_Product12_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1110_out;
SharedReg86_out_to_MUX_Product12_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg86_out;
SharedReg1146_out_to_MUX_Product12_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1146_out;
SharedReg1104_out_to_MUX_Product12_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1104_out;
SharedReg1133_out_to_MUX_Product12_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1133_out;
SharedReg1151_out_to_MUX_Product12_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1151_out;
SharedReg86_out_to_MUX_Product12_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg86_out;
SharedReg89_out_to_MUX_Product12_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg89_out;
SharedReg286_out_to_MUX_Product12_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg286_out;
SharedReg183_out_to_MUX_Product12_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg183_out;
SharedReg182_out_to_MUX_Product12_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg182_out;
   MUX_Product12_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg118_out_to_MUX_Product12_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1110_out_to_MUX_Product12_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg183_out_to_MUX_Product12_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg182_out_to_MUX_Product12_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg86_out_to_MUX_Product12_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1146_out_to_MUX_Product12_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1104_out_to_MUX_Product12_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1133_out_to_MUX_Product12_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1151_out_to_MUX_Product12_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg86_out_to_MUX_Product12_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg89_out_to_MUX_Product12_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg286_out_to_MUX_Product12_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product12_5_impl_0_out);

   Delay1No230_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_5_impl_0_out,
                 Y => Delay1No230_out);

SharedReg1124_out_to_MUX_Product12_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1124_out;
SharedReg89_out_to_MUX_Product12_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg89_out;
SharedReg1126_out_to_MUX_Product12_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1126_out;
SharedReg1060_out_to_MUX_Product12_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1060_out;
SharedReg151_out_to_MUX_Product12_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg151_out;
SharedReg999_out_to_MUX_Product12_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg999_out;
SharedReg1061_out_to_MUX_Product12_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1061_out;
SharedReg1119_out_to_MUX_Product12_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product12_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1125_out;
SharedReg1120_out_to_MUX_Product12_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1120_out;
SharedReg1121_out_to_MUX_Product12_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1121_out;
SharedReg1123_out_to_MUX_Product12_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1123_out;
   MUX_Product12_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1124_out_to_MUX_Product12_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg89_out_to_MUX_Product12_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1121_out_to_MUX_Product12_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1123_out_to_MUX_Product12_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1126_out_to_MUX_Product12_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1060_out_to_MUX_Product12_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg151_out_to_MUX_Product12_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg999_out_to_MUX_Product12_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1061_out_to_MUX_Product12_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1119_out_to_MUX_Product12_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1125_out_to_MUX_Product12_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1120_out_to_MUX_Product12_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product12_5_impl_1_out);

   Delay1No231_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_5_impl_1_out,
                 Y => Delay1No231_out);

Delay1No232_out_to_Product12_6_impl_parent_implementedSystem_port_0_cast <= Delay1No232_out;
Delay1No233_out_to_Product12_6_impl_parent_implementedSystem_port_1_cast <= Delay1No233_out;
   Product12_6_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product12_6_impl_out,
                 X => Delay1No232_out_to_Product12_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No233_out_to_Product12_6_impl_parent_implementedSystem_port_1_cast);

SharedReg123_out_to_MUX_Product12_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg123_out;
SharedReg123_out_to_MUX_Product12_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg123_out;
SharedReg1110_out_to_MUX_Product12_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1110_out;
SharedReg60_out_to_MUX_Product12_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg60_out;
SharedReg1146_out_to_MUX_Product12_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1146_out;
SharedReg1104_out_to_MUX_Product12_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1104_out;
SharedReg1133_out_to_MUX_Product12_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1133_out;
SharedReg1151_out_to_MUX_Product12_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1151_out;
SharedReg91_out_to_MUX_Product12_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg91_out;
SharedReg125_out_to_MUX_Product12_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg125_out;
SharedReg218_out_to_MUX_Product12_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg218_out;
SharedReg154_out_to_MUX_Product12_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg154_out;
   MUX_Product12_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg123_out_to_MUX_Product12_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg123_out_to_MUX_Product12_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg218_out_to_MUX_Product12_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg154_out_to_MUX_Product12_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1110_out_to_MUX_Product12_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg60_out_to_MUX_Product12_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1146_out_to_MUX_Product12_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1104_out_to_MUX_Product12_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1133_out_to_MUX_Product12_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1151_out_to_MUX_Product12_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg91_out_to_MUX_Product12_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg125_out_to_MUX_Product12_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product12_6_impl_0_out);

   Delay1No232_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_6_impl_0_out,
                 Y => Delay1No232_out);

SharedReg1123_out_to_MUX_Product12_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1123_out;
SharedReg1124_out_to_MUX_Product12_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1124_out;
SharedReg94_out_to_MUX_Product12_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg94_out;
SharedReg1126_out_to_MUX_Product12_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1126_out;
SharedReg1088_out_to_MUX_Product12_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1088_out;
SharedReg154_out_to_MUX_Product12_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg154_out;
SharedReg1068_out_to_MUX_Product12_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1068_out;
SharedReg1077_out_to_MUX_Product12_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1077_out;
SharedReg1119_out_to_MUX_Product12_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product12_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1125_out;
SharedReg1120_out_to_MUX_Product12_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1120_out;
SharedReg1121_out_to_MUX_Product12_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1121_out;
   MUX_Product12_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1123_out_to_MUX_Product12_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1124_out_to_MUX_Product12_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1120_out_to_MUX_Product12_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1121_out_to_MUX_Product12_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg94_out_to_MUX_Product12_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1126_out_to_MUX_Product12_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1088_out_to_MUX_Product12_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg154_out_to_MUX_Product12_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1068_out_to_MUX_Product12_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1077_out_to_MUX_Product12_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1119_out_to_MUX_Product12_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1125_out_to_MUX_Product12_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product12_6_impl_1_out);

   Delay1No233_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_6_impl_1_out,
                 Y => Delay1No233_out);

Delay1No234_out_to_Product22_0_impl_parent_implementedSystem_port_0_cast <= Delay1No234_out;
Delay1No235_out_to_Product22_0_impl_parent_implementedSystem_port_1_cast <= Delay1No235_out;
   Product22_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product22_0_impl_out,
                 X => Delay1No234_out_to_Product22_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No235_out_to_Product22_0_impl_parent_implementedSystem_port_1_cast);

SharedReg1108_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1108_out;
SharedReg1109_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1109_out;
SharedReg1136_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1136_out;
SharedReg1112_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1112_out;
SharedReg1122_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1122_out;
SharedReg1114_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1114_out;
SharedReg1094_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1094_out;
SharedReg1116_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1116_out;
SharedReg1134_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1134_out;
SharedReg1106_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1106_out;
SharedReg1107_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1113_out;
   MUX_Product22_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1108_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1109_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1107_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1113_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1136_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1112_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1122_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1114_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1094_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1116_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1134_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1106_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product22_0_impl_0_out);

   Delay1No234_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product22_0_impl_0_out,
                 Y => Delay1No234_out);

SharedReg65_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg65_out;
SharedReg33_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg33_out;
SharedReg564_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg564_out;
SharedReg95_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg95_out;
SharedReg204_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg204_out;
SharedReg205_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg205_out;
SharedReg1150_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1150_out;
SharedReg96_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg96_out;
SharedReg1005_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1005_out;
SharedReg67_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg67_out;
SharedReg95_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg95_out;
SharedReg35_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg35_out;
   MUX_Product22_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg65_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg33_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg95_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg35_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg564_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg95_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg204_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg205_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1150_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg96_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1005_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg67_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product22_0_impl_1_out);

   Delay1No235_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product22_0_impl_1_out,
                 Y => Delay1No235_out);

Delay1No236_out_to_Product22_1_impl_parent_implementedSystem_port_0_cast <= Delay1No236_out;
Delay1No237_out_to_Product22_1_impl_parent_implementedSystem_port_1_cast <= Delay1No237_out;
   Product22_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product22_1_impl_out,
                 X => Delay1No236_out_to_Product22_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No237_out_to_Product22_1_impl_parent_implementedSystem_port_1_cast);

SharedReg1107_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1113_out;
SharedReg1108_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1108_out;
SharedReg1109_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1109_out;
SharedReg1136_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1136_out;
SharedReg1112_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1112_out;
SharedReg1122_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1122_out;
SharedReg1114_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1114_out;
SharedReg783_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg783_out;
SharedReg1116_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1116_out;
SharedReg1134_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1134_out;
SharedReg1106_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1106_out;
   MUX_Product22_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1107_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1113_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1134_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1106_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1108_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1109_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1136_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1112_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1122_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1114_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg783_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1116_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product22_1_impl_0_out);

   Delay1No236_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product22_1_impl_0_out,
                 Y => Delay1No236_out);

SharedReg69_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg69_out;
SharedReg161_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg161_out;
SharedReg38_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg38_out;
SharedReg159_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg159_out;
SharedReg438_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg438_out;
SharedReg69_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg69_out;
SharedReg132_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg132_out;
SharedReg133_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg133_out;
SharedReg1150_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1150_out;
SharedReg101_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg101_out;
SharedReg1008_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1008_out;
SharedReg71_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg71_out;
   MUX_Product22_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg69_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg161_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1008_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg71_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg38_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg159_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg438_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg69_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg132_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg133_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1150_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg101_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product22_1_impl_1_out);

   Delay1No237_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product22_1_impl_1_out,
                 Y => Delay1No237_out);

Delay1No238_out_to_Product22_2_impl_parent_implementedSystem_port_0_cast <= Delay1No238_out;
Delay1No239_out_to_Product22_2_impl_parent_implementedSystem_port_1_cast <= Delay1No239_out;
   Product22_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product22_2_impl_out,
                 X => Delay1No238_out_to_Product22_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No239_out_to_Product22_2_impl_parent_implementedSystem_port_1_cast);

SharedReg1134_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1134_out;
SharedReg1106_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1106_out;
SharedReg1107_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1113_out;
SharedReg1108_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1108_out;
SharedReg1109_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1109_out;
SharedReg1136_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1136_out;
SharedReg1112_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1112_out;
SharedReg1122_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1122_out;
SharedReg1114_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1114_out;
SharedReg876_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg876_out;
SharedReg1116_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1116_out;
   MUX_Product22_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1134_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1106_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg876_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1116_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1107_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1113_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1108_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1109_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1136_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1112_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1122_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1114_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product22_2_impl_0_out);

   Delay1No238_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product22_2_impl_0_out,
                 Y => Delay1No238_out);

SharedReg987_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg987_out;
SharedReg75_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg75_out;
SharedReg73_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg73_out;
SharedReg166_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg166_out;
SharedReg41_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg41_out;
SharedReg165_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg165_out;
SharedReg445_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg445_out;
SharedReg105_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg105_out;
SharedReg136_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg136_out;
SharedReg138_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg138_out;
SharedReg1150_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1150_out;
SharedReg106_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg106_out;
   MUX_Product22_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg987_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg75_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1150_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg106_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg73_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg166_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg41_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg165_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg445_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg105_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg136_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg138_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product22_2_impl_1_out);

   Delay1No239_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product22_2_impl_1_out,
                 Y => Delay1No239_out);

Delay1No240_out_to_Product22_3_impl_parent_implementedSystem_port_0_cast <= Delay1No240_out;
Delay1No241_out_to_Product22_3_impl_parent_implementedSystem_port_1_cast <= Delay1No241_out;
   Product22_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product22_3_impl_out,
                 X => Delay1No240_out_to_Product22_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No241_out_to_Product22_3_impl_parent_implementedSystem_port_1_cast);

SharedReg1116_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1116_out;
SharedReg1134_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1134_out;
SharedReg1106_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1106_out;
SharedReg1107_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1113_out;
SharedReg1108_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1108_out;
SharedReg1109_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1109_out;
SharedReg1136_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1136_out;
SharedReg1112_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1112_out;
SharedReg1122_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1122_out;
SharedReg1114_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1114_out;
SharedReg758_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg758_out;
   MUX_Product22_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1116_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1134_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1114_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg758_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1106_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1107_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1113_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1108_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1109_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1136_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1112_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1122_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product22_3_impl_0_out);

   Delay1No240_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product22_3_impl_0_out,
                 Y => Delay1No240_out);

SharedReg111_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg111_out;
SharedReg991_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg991_out;
SharedReg46_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg46_out;
SharedReg44_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg44_out;
SharedReg200_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg200_out;
SharedReg198_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg198_out;
SharedReg171_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg171_out;
SharedReg451_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg451_out;
SharedReg110_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg110_out;
SharedReg142_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg142_out;
SharedReg113_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg113_out;
SharedReg1150_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1150_out;
   MUX_Product22_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg111_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg991_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg113_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1150_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg46_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg44_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg200_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg198_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg171_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg451_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg110_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg142_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product22_3_impl_1_out);

   Delay1No241_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product22_3_impl_1_out,
                 Y => Delay1No241_out);

Delay1No242_out_to_Product22_4_impl_parent_implementedSystem_port_0_cast <= Delay1No242_out;
Delay1No243_out_to_Product22_4_impl_parent_implementedSystem_port_1_cast <= Delay1No243_out;
   Product22_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product22_4_impl_out,
                 X => Delay1No242_out_to_Product22_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No243_out_to_Product22_4_impl_parent_implementedSystem_port_1_cast);

SharedReg1114_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1114_out;
SharedReg764_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg764_out;
SharedReg1116_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1116_out;
SharedReg1134_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1134_out;
SharedReg1106_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1106_out;
SharedReg1107_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1113_out;
SharedReg1108_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1108_out;
SharedReg1109_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1109_out;
SharedReg1136_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1136_out;
SharedReg1112_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1112_out;
SharedReg1122_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1122_out;
   MUX_Product22_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1114_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg764_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1112_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1122_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1116_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1134_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1106_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1107_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1113_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1108_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1109_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1136_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product22_4_impl_0_out);

   Delay1No242_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product22_4_impl_0_out,
                 Y => Delay1No242_out);

SharedReg117_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg117_out;
SharedReg1150_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1150_out;
SharedReg115_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg115_out;
SharedReg866_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg866_out;
SharedReg50_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg50_out;
SharedReg48_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg48_out;
SharedReg193_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg193_out;
SharedReg48_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg48_out;
SharedReg176_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg176_out;
SharedReg458_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg458_out;
SharedReg114_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg114_out;
SharedReg209_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg209_out;
   MUX_Product22_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg117_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1150_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg114_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg209_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg115_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg866_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg50_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg48_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg193_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg48_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg176_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg458_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product22_4_impl_1_out);

   Delay1No243_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product22_4_impl_1_out,
                 Y => Delay1No243_out);

Delay1No244_out_to_Product22_5_impl_parent_implementedSystem_port_0_cast <= Delay1No244_out;
Delay1No245_out_to_Product22_5_impl_parent_implementedSystem_port_1_cast <= Delay1No245_out;
   Product22_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product22_5_impl_out,
                 X => Delay1No244_out_to_Product22_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No245_out_to_Product22_5_impl_parent_implementedSystem_port_1_cast);

SharedReg1112_out_to_MUX_Product22_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1112_out;
SharedReg1122_out_to_MUX_Product22_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1122_out;
SharedReg1114_out_to_MUX_Product22_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1114_out;
SharedReg1060_out_to_MUX_Product22_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1060_out;
SharedReg1116_out_to_MUX_Product22_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1116_out;
SharedReg1134_out_to_MUX_Product22_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1134_out;
SharedReg1106_out_to_MUX_Product22_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1106_out;
SharedReg1107_out_to_MUX_Product22_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product22_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1113_out;
SharedReg1108_out_to_MUX_Product22_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1108_out;
SharedReg1109_out_to_MUX_Product22_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1109_out;
SharedReg1136_out_to_MUX_Product22_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1136_out;
   MUX_Product22_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1112_out_to_MUX_Product22_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1122_out_to_MUX_Product22_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1109_out_to_MUX_Product22_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1136_out_to_MUX_Product22_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1114_out_to_MUX_Product22_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1060_out_to_MUX_Product22_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1116_out_to_MUX_Product22_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1134_out_to_MUX_Product22_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1106_out_to_MUX_Product22_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1107_out_to_MUX_Product22_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1113_out_to_MUX_Product22_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1108_out_to_MUX_Product22_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product22_5_impl_0_out);

   Delay1No244_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product22_5_impl_0_out,
                 Y => Delay1No244_out);

SharedReg150_out_to_MUX_Product22_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg150_out;
SharedReg215_out_to_MUX_Product22_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg215_out;
SharedReg186_out_to_MUX_Product22_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg186_out;
SharedReg1150_out_to_MUX_Product22_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1150_out;
SharedReg119_out_to_MUX_Product22_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg119_out;
SharedReg869_out_to_MUX_Product22_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg869_out;
SharedReg88_out_to_MUX_Product22_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg88_out;
SharedReg118_out_to_MUX_Product22_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg118_out;
SharedReg281_out_to_MUX_Product22_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg281_out;
SharedReg118_out_to_MUX_Product22_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg118_out;
SharedReg87_out_to_MUX_Product22_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg87_out;
SharedReg589_out_to_MUX_Product22_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg589_out;
   MUX_Product22_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg150_out_to_MUX_Product22_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg215_out_to_MUX_Product22_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg87_out_to_MUX_Product22_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg589_out_to_MUX_Product22_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg186_out_to_MUX_Product22_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1150_out_to_MUX_Product22_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg119_out_to_MUX_Product22_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg869_out_to_MUX_Product22_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg88_out_to_MUX_Product22_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg118_out_to_MUX_Product22_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg281_out_to_MUX_Product22_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg118_out_to_MUX_Product22_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product22_5_impl_1_out);

   Delay1No245_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product22_5_impl_1_out,
                 Y => Delay1No245_out);

Delay1No246_out_to_Product22_6_impl_parent_implementedSystem_port_0_cast <= Delay1No246_out;
Delay1No247_out_to_Product22_6_impl_parent_implementedSystem_port_1_cast <= Delay1No247_out;
   Product22_6_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product22_6_impl_out,
                 X => Delay1No246_out_to_Product22_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No247_out_to_Product22_6_impl_parent_implementedSystem_port_1_cast);

SharedReg1136_out_to_MUX_Product22_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1136_out;
SharedReg1112_out_to_MUX_Product22_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1112_out;
SharedReg1122_out_to_MUX_Product22_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1122_out;
SharedReg1114_out_to_MUX_Product22_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1114_out;
SharedReg1088_out_to_MUX_Product22_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1088_out;
SharedReg1116_out_to_MUX_Product22_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1116_out;
SharedReg1134_out_to_MUX_Product22_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1134_out;
SharedReg1106_out_to_MUX_Product22_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1106_out;
SharedReg1107_out_to_MUX_Product22_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product22_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1113_out;
SharedReg1108_out_to_MUX_Product22_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1108_out;
SharedReg1109_out_to_MUX_Product22_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1109_out;
   MUX_Product22_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1136_out_to_MUX_Product22_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1112_out_to_MUX_Product22_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1108_out_to_MUX_Product22_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1109_out_to_MUX_Product22_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1122_out_to_MUX_Product22_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1114_out_to_MUX_Product22_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1088_out_to_MUX_Product22_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1116_out_to_MUX_Product22_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1134_out_to_MUX_Product22_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1106_out_to_MUX_Product22_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1107_out_to_MUX_Product22_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1113_out_to_MUX_Product22_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product22_6_impl_0_out);

   Delay1No246_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product22_6_impl_0_out,
                 Y => Delay1No246_out);

SharedReg595_out_to_MUX_Product22_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg595_out;
SharedReg153_out_to_MUX_Product22_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg153_out;
SharedReg221_out_to_MUX_Product22_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg221_out;
SharedReg190_out_to_MUX_Product22_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg190_out;
SharedReg1150_out_to_MUX_Product22_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1150_out;
SharedReg124_out_to_MUX_Product22_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg124_out;
SharedReg1002_out_to_MUX_Product22_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1002_out;
SharedReg62_out_to_MUX_Product22_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg62_out;
SharedReg123_out_to_MUX_Product22_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg123_out;
SharedReg63_out_to_MUX_Product22_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg63_out;
SharedReg91_out_to_MUX_Product22_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg91_out;
SharedReg61_out_to_MUX_Product22_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg61_out;
   MUX_Product22_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg595_out_to_MUX_Product22_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg153_out_to_MUX_Product22_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg91_out_to_MUX_Product22_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg61_out_to_MUX_Product22_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg221_out_to_MUX_Product22_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg190_out_to_MUX_Product22_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1150_out_to_MUX_Product22_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg124_out_to_MUX_Product22_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1002_out_to_MUX_Product22_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg62_out_to_MUX_Product22_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg123_out_to_MUX_Product22_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg63_out_to_MUX_Product22_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product22_6_impl_1_out);

   Delay1No247_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product22_6_impl_1_out,
                 Y => Delay1No247_out);

Delay1No248_out_to_Product32_0_impl_parent_implementedSystem_port_0_cast <= Delay1No248_out;
Delay1No249_out_to_Product32_0_impl_parent_implementedSystem_port_1_cast <= Delay1No249_out;
   Product32_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_0_impl_out,
                 X => Delay1No248_out_to_Product32_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No249_out_to_Product32_0_impl_parent_implementedSystem_port_1_cast);

SharedReg1108_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1108_out;
SharedReg1109_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1109_out;
SharedReg1136_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1136_out;
SharedReg1112_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1112_out;
SharedReg35_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg35_out;
SharedReg1114_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1114_out;
SharedReg1154_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1154_out;
SharedReg128_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg128_out;
SharedReg1134_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1134_out;
SharedReg67_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg67_out;
SharedReg1107_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1113_out;
   MUX_Product32_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1108_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1109_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1107_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1113_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1136_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1112_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg35_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1114_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1154_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg128_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1134_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg67_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product32_0_impl_0_out);

   Delay1No248_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_0_impl_0_out,
                 Y => Delay1No248_out);

SharedReg95_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg95_out;
SharedReg127_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg127_out;
SharedReg666_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg666_out;
SharedReg127_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg127_out;
SharedReg1122_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1122_out;
SharedReg36_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg36_out;
SharedReg775_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg775_out;
SharedReg1116_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1116_out;
SharedReg1038_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1038_out;
SharedReg1118_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1118_out;
SharedReg127_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg127_out;
SharedReg68_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg68_out;
   MUX_Product32_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg95_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg127_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg127_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg68_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg666_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg127_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1122_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg36_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg775_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1116_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1038_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1118_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product32_0_impl_1_out);

   Delay1No249_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_0_impl_1_out,
                 Y => Delay1No249_out);

Delay1No250_out_to_Product32_1_impl_parent_implementedSystem_port_0_cast <= Delay1No250_out;
Delay1No251_out_to_Product32_1_impl_parent_implementedSystem_port_1_cast <= Delay1No251_out;
   Product32_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_1_impl_out,
                 X => Delay1No250_out_to_Product32_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No251_out_to_Product32_1_impl_parent_implementedSystem_port_1_cast);

SharedReg1107_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1113_out;
SharedReg1108_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1108_out;
SharedReg1109_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1109_out;
SharedReg1136_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1136_out;
SharedReg1112_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1112_out;
SharedReg161_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg161_out;
SharedReg1114_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1114_out;
SharedReg1154_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1154_out;
SharedReg131_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg131_out;
SharedReg1134_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1134_out;
SharedReg71_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg71_out;
   MUX_Product32_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1107_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1113_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1134_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg71_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1108_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1109_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1136_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1112_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg161_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1114_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1154_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg131_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product32_1_impl_0_out);

   Delay1No250_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_1_impl_0_out,
                 Y => Delay1No250_out);

SharedReg100_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg100_out;
SharedReg40_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg40_out;
SharedReg69_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg69_out;
SharedReg100_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg100_out;
SharedReg570_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg570_out;
SharedReg100_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg100_out;
SharedReg1122_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1122_out;
SharedReg162_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg162_out;
SharedReg746_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg746_out;
SharedReg1116_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1116_out;
SharedReg1043_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1043_out;
SharedReg1118_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1118_out;
   MUX_Product32_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg100_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg40_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1043_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1118_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg69_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg100_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg570_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg100_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1122_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg162_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg746_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1116_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product32_1_impl_1_out);

   Delay1No251_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_1_impl_1_out,
                 Y => Delay1No251_out);

Delay1No252_out_to_Product32_2_impl_parent_implementedSystem_port_0_cast <= Delay1No252_out;
Delay1No253_out_to_Product32_2_impl_parent_implementedSystem_port_1_cast <= Delay1No253_out;
   Product32_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_2_impl_out,
                 X => Delay1No252_out_to_Product32_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No253_out_to_Product32_2_impl_parent_implementedSystem_port_1_cast);

SharedReg1134_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1134_out;
SharedReg75_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg75_out;
SharedReg1107_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1113_out;
SharedReg1108_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1108_out;
SharedReg1109_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1109_out;
SharedReg1136_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1136_out;
SharedReg1112_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1112_out;
SharedReg166_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg166_out;
SharedReg1114_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1114_out;
SharedReg1154_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1154_out;
SharedReg135_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg135_out;
   MUX_Product32_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1134_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg75_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1154_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg135_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1107_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1113_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1108_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1109_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1136_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1112_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg166_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1114_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product32_2_impl_0_out);

   Delay1No252_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_2_impl_0_out,
                 Y => Delay1No252_out);

SharedReg1013_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1013_out;
SharedReg1118_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1118_out;
SharedReg105_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg105_out;
SharedReg43_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg43_out;
SharedReg73_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg73_out;
SharedReg105_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg105_out;
SharedReg576_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg576_out;
SharedReg134_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg134_out;
SharedReg1122_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1122_out;
SharedReg167_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg167_out;
SharedReg753_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg753_out;
SharedReg1116_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1116_out;
   MUX_Product32_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1013_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1118_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg753_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1116_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg105_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg43_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg73_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg105_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg576_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg134_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1122_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg167_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product32_2_impl_1_out);

   Delay1No253_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_2_impl_1_out,
                 Y => Delay1No253_out);

Delay1No254_out_to_Product32_3_impl_parent_implementedSystem_port_0_cast <= Delay1No254_out;
Delay1No255_out_to_Product32_3_impl_parent_implementedSystem_port_1_cast <= Delay1No255_out;
   Product32_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_3_impl_out,
                 X => Delay1No254_out_to_Product32_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No255_out_to_Product32_3_impl_parent_implementedSystem_port_1_cast);

SharedReg140_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg140_out;
SharedReg1134_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1134_out;
SharedReg46_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg46_out;
SharedReg1107_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1113_out;
SharedReg1108_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1108_out;
SharedReg1109_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1109_out;
SharedReg1136_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1136_out;
SharedReg1112_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1112_out;
SharedReg200_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg200_out;
SharedReg1114_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1114_out;
SharedReg1154_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1154_out;
   MUX_Product32_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg140_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1134_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1114_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1154_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg46_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1107_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1113_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1108_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1109_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1136_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1112_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg200_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product32_3_impl_0_out);

   Delay1No254_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_3_impl_0_out,
                 Y => Delay1No254_out);

SharedReg1116_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1116_out;
SharedReg1018_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1018_out;
SharedReg1118_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1118_out;
SharedReg77_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg77_out;
SharedReg47_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg47_out;
SharedReg44_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg44_out;
SharedReg110_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg110_out;
SharedReg580_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg580_out;
SharedReg139_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg139_out;
SharedReg1122_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1122_out;
SharedReg172_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg172_out;
SharedReg705_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg705_out;
   MUX_Product32_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1116_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1018_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg172_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg705_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1118_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg77_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg47_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg44_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg110_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg580_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg139_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1122_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product32_3_impl_1_out);

   Delay1No255_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_3_impl_1_out,
                 Y => Delay1No255_out);

Delay1No256_out_to_Product32_4_impl_parent_implementedSystem_port_0_cast <= Delay1No256_out;
Delay1No257_out_to_Product32_4_impl_parent_implementedSystem_port_1_cast <= Delay1No257_out;
   Product32_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_4_impl_out,
                 X => Delay1No256_out_to_Product32_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No257_out_to_Product32_4_impl_parent_implementedSystem_port_1_cast);

SharedReg1114_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1114_out;
SharedReg1154_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1154_out;
SharedReg146_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg146_out;
SharedReg1134_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1134_out;
SharedReg50_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg50_out;
SharedReg1107_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1113_out;
SharedReg1108_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1108_out;
SharedReg1109_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1109_out;
SharedReg1136_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1136_out;
SharedReg1112_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1112_out;
SharedReg51_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg51_out;
   MUX_Product32_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1114_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1154_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1112_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg51_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg146_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1134_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg50_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1107_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1113_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1108_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1109_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1136_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product32_4_impl_0_out);

   Delay1No256_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_4_impl_0_out,
                 Y => Delay1No256_out);

SharedReg179_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg179_out;
SharedReg712_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg712_out;
SharedReg1116_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1116_out;
SharedReg994_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg994_out;
SharedReg1118_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1118_out;
SharedReg81_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg81_out;
SharedReg178_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg178_out;
SharedReg81_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg81_out;
SharedReg145_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg145_out;
SharedReg584_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg584_out;
SharedReg145_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg145_out;
SharedReg1122_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1122_out;
   MUX_Product32_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg179_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg712_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg145_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1122_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1116_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg994_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1118_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg81_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg178_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg81_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg145_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg584_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product32_4_impl_1_out);

   Delay1No257_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_4_impl_1_out,
                 Y => Delay1No257_out);

Delay1No258_out_to_Product32_5_impl_parent_implementedSystem_port_0_cast <= Delay1No258_out;
Delay1No259_out_to_Product32_5_impl_parent_implementedSystem_port_1_cast <= Delay1No259_out;
   Product32_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_5_impl_out,
                 X => Delay1No258_out_to_Product32_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No259_out_to_Product32_5_impl_parent_implementedSystem_port_1_cast);

SharedReg1112_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1112_out;
SharedReg89_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg89_out;
SharedReg1114_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1114_out;
SharedReg1154_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1154_out;
SharedReg151_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg151_out;
SharedReg1134_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1134_out;
SharedReg88_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg88_out;
SharedReg1107_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1113_out;
SharedReg1108_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1108_out;
SharedReg1109_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1109_out;
SharedReg1136_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1136_out;
   MUX_Product32_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1112_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg89_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1109_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1136_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1114_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1154_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg151_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1134_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg88_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1107_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1113_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1108_out_to_MUX_Product32_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product32_5_impl_0_out);

   Delay1No258_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_5_impl_0_out,
                 Y => Delay1No258_out);

SharedReg182_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg182_out;
SharedReg1122_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1122_out;
SharedReg90_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg90_out;
SharedReg770_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg770_out;
SharedReg1116_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1116_out;
SharedReg998_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg998_out;
SharedReg1118_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1118_out;
SharedReg150_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg150_out;
SharedReg55_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg55_out;
SharedReg150_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg150_out;
SharedReg182_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg182_out;
SharedReg694_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg694_out;
   MUX_Product32_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg182_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1122_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg182_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg694_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg90_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg770_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1116_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg998_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1118_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg150_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg55_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg150_out_to_MUX_Product32_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product32_5_impl_1_out);

   Delay1No259_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_5_impl_1_out,
                 Y => Delay1No259_out);

Delay1No260_out_to_Product32_6_impl_parent_implementedSystem_port_0_cast <= Delay1No260_out;
Delay1No261_out_to_Product32_6_impl_parent_implementedSystem_port_1_cast <= Delay1No261_out;
   Product32_6_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_6_impl_out,
                 X => Delay1No260_out_to_Product32_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No261_out_to_Product32_6_impl_parent_implementedSystem_port_1_cast);

SharedReg1136_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1136_out;
SharedReg1112_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1112_out;
SharedReg94_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg94_out;
SharedReg1114_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1114_out;
SharedReg1154_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1154_out;
SharedReg154_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg154_out;
SharedReg1134_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1134_out;
SharedReg62_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg62_out;
SharedReg1107_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1113_out;
SharedReg1108_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1108_out;
SharedReg1109_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1109_out;
   MUX_Product32_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1136_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1112_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1108_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1109_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg94_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1114_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1154_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg154_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1134_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg62_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1107_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1113_out_to_MUX_Product32_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product32_6_impl_0_out);

   Delay1No260_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_6_impl_0_out,
                 Y => Delay1No260_out);

SharedReg699_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg699_out;
SharedReg187_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg187_out;
SharedReg1122_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1122_out;
SharedReg64_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg64_out;
SharedReg1101_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1101_out;
SharedReg1116_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1116_out;
SharedReg1034_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1034_out;
SharedReg1118_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1118_out;
SharedReg153_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg153_out;
SharedReg94_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg94_out;
SharedReg123_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg123_out;
SharedReg187_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg187_out;
   MUX_Product32_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg699_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg187_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg123_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg187_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1122_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg64_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1101_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1116_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1034_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1118_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg153_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg94_out_to_MUX_Product32_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product32_6_impl_1_out);

   Delay1No261_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_6_impl_1_out,
                 Y => Delay1No261_out);

Delay1No262_out_to_Subtract3_0_impl_parent_implementedSystem_port_0_cast <= Delay1No262_out;
Delay1No263_out_to_Subtract3_0_impl_parent_implementedSystem_port_1_cast <= Delay1No263_out;
   Subtract3_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract3_0_impl_out,
                 X => Delay1No262_out_to_Subtract3_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No263_out_to_Subtract3_0_impl_parent_implementedSystem_port_1_cast);

SharedReg529_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg529_out;
SharedReg1_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1_out;
SharedReg720_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg720_out;
SharedReg396_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg396_out;
SharedReg529_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg529_out;
SharedReg529_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg529_out;
SharedReg529_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg529_out;
SharedReg529_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg529_out;
SharedReg883_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg883_out;
SharedReg564_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg564_out;
SharedReg431_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg431_out;
SharedReg480_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg480_out;
   MUX_Subtract3_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg529_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg431_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg480_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg720_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg396_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg529_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg529_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg529_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg529_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg883_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg564_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract3_0_impl_0_out);

   Delay1No262_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_0_impl_0_out,
                 Y => Delay1No262_out);

SharedReg624_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg624_out;
SharedReg17_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg17_out;
SharedReg551_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg551_out;
SharedReg502_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg502_out;
SharedReg624_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg624_out;
SharedReg624_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg624_out;
SharedReg624_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg624_out;
SharedReg624_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg624_out;
SharedReg960_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg960_out;
SharedReg667_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg667_out;
SharedReg564_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg564_out;
SharedReg550_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg550_out;
   MUX_Subtract3_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg624_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg17_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg564_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg550_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg551_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg502_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg624_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg624_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg624_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg624_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg960_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg667_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract3_0_impl_1_out);

   Delay1No263_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_0_impl_1_out,
                 Y => Delay1No263_out);

Delay1No264_out_to_Subtract3_1_impl_parent_implementedSystem_port_0_cast <= Delay1No264_out;
Delay1No265_out_to_Subtract3_1_impl_parent_implementedSystem_port_1_cast <= Delay1No265_out;
   Subtract3_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract3_1_impl_out,
                 X => Delay1No264_out_to_Subtract3_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No265_out_to_Subtract3_1_impl_parent_implementedSystem_port_1_cast);

SharedReg70_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg70_out;
SharedReg483_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg483_out;
SharedReg532_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg532_out;
SharedReg1_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1_out;
SharedReg724_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg724_out;
SharedReg533_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg533_out;
SharedReg648_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg648_out;
SharedReg648_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg648_out;
SharedReg1009_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1009_out;
SharedReg648_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg648_out;
SharedReg888_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg888_out;
SharedReg100_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg100_out;
   MUX_Subtract3_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg70_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg483_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg888_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg100_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg532_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg724_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg533_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg648_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg648_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1009_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg648_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract3_1_impl_0_out);

   Delay1No264_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_1_impl_0_out,
                 Y => Delay1No264_out);

SharedReg254_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg254_out;
SharedReg552_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg552_out;
SharedReg627_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg627_out;
SharedReg17_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg17_out;
SharedReg553_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg553_out;
SharedReg628_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg628_out;
SharedReg825_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg825_out;
SharedReg825_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg825_out;
SharedReg444_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg444_out;
SharedReg825_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg825_out;
SharedReg964_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg964_out;
SharedReg235_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg235_out;
   MUX_Subtract3_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg254_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg552_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg964_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg235_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg627_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg17_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg553_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg628_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg825_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg825_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg444_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg825_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract3_1_impl_1_out);

   Delay1No265_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_1_impl_1_out,
                 Y => Delay1No265_out);

Delay1No266_out_to_Subtract3_2_impl_parent_implementedSystem_port_0_cast <= Delay1No266_out;
Delay1No267_out_to_Subtract3_2_impl_parent_implementedSystem_port_1_cast <= Delay1No267_out;
   Subtract3_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract3_2_impl_out,
                 X => Delay1No266_out_to_Subtract3_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No267_out_to_Subtract3_2_impl_parent_implementedSystem_port_1_cast);

SharedReg749_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg749_out;
SharedReg105_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg105_out;
SharedReg74_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg74_out;
SharedReg486_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg486_out;
SharedReg535_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg535_out;
SharedReg2_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg2_out;
SharedReg652_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg652_out;
SharedReg652_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg652_out;
SharedReg891_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg891_out;
SharedReg891_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg891_out;
SharedReg304_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg304_out;
SharedReg445_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg445_out;
   MUX_Subtract3_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg749_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg105_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg304_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg445_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg74_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg486_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg535_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg2_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg652_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg652_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg891_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg891_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract3_2_impl_0_out);

   Delay1No266_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_2_impl_0_out,
                 Y => Delay1No266_out);

SharedReg986_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg986_out;
SharedReg240_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg240_out;
SharedReg260_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg260_out;
SharedReg554_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg554_out;
SharedReg630_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg630_out;
SharedReg18_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg18_out;
SharedReg830_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg830_out;
SharedReg830_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg830_out;
SharedReg966_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg966_out;
SharedReg966_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg966_out;
SharedReg307_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg307_out;
SharedReg678_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg678_out;
   MUX_Subtract3_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg986_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg240_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg307_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg678_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg260_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg554_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg630_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg18_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg830_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg830_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg966_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg966_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract3_2_impl_1_out);

   Delay1No267_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_2_impl_1_out,
                 Y => Delay1No267_out);

Delay1No268_out_to_Subtract3_3_impl_parent_implementedSystem_port_0_cast <= Delay1No268_out;
Delay1No269_out_to_Subtract3_3_impl_parent_implementedSystem_port_1_cast <= Delay1No269_out;
   Subtract3_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract3_3_impl_out,
                 X => Delay1No268_out_to_Subtract3_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No269_out_to_Subtract3_3_impl_parent_implementedSystem_port_1_cast);

SharedReg451_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg451_out;
SharedReg896_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg896_out;
SharedReg77_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg77_out;
SharedReg877_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg877_out;
SharedReg489_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg489_out;
SharedReg538_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg538_out;
SharedReg1_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1_out;
SharedReg655_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg655_out;
SharedReg539_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg539_out;
SharedReg895_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg895_out;
SharedReg895_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg895_out;
SharedReg267_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg267_out;
   MUX_Subtract3_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg451_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg896_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg895_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg267_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg77_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg877_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg489_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg538_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg655_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg539_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg895_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract3_3_impl_0_out);

   Delay1No268_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_3_impl_0_out,
                 Y => Delay1No268_out);

SharedReg683_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg683_out;
SharedReg970_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg970_out;
SharedReg245_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg245_out;
SharedReg753_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg753_out;
SharedReg556_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg556_out;
SharedReg633_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg633_out;
SharedReg17_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg17_out;
SharedReg834_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg834_out;
SharedReg634_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg634_out;
SharedReg969_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg969_out;
SharedReg969_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg969_out;
SharedReg271_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg271_out;
   MUX_Subtract3_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg683_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg970_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg969_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg271_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg245_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg753_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg556_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg633_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg17_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg834_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg634_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg969_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract3_3_impl_1_out);

   Delay1No269_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_3_impl_1_out,
                 Y => Delay1No269_out);

Delay1No270_out_to_Subtract3_4_impl_parent_implementedSystem_port_0_cast <= Delay1No270_out;
Delay1No271_out_to_Subtract3_4_impl_parent_implementedSystem_port_1_cast <= Delay1No271_out;
   Subtract3_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract3_4_impl_out,
                 X => Delay1No270_out_to_Subtract3_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No271_out_to_Subtract3_4_impl_parent_implementedSystem_port_1_cast);

SharedReg993_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg993_out;
SharedReg310_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg310_out;
SharedReg705_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg705_out;
SharedReg900_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg900_out;
SharedReg81_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg81_out;
SharedReg49_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg49_out;
SharedReg492_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg492_out;
Delay4No214_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_8_cast <= Delay4No214_out;
SharedReg2_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg2_out;
SharedReg952_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg952_out;
SharedReg900_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg900_out;
SharedReg542_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg542_out;
   MUX_Subtract3_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg993_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg310_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg900_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg542_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg705_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg900_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg81_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg49_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg492_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay4No214_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg2_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg952_out_to_MUX_Subtract3_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract3_4_impl_0_out);

   Delay1No270_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_4_impl_0_out,
                 Y => Delay1No270_out);

SharedReg458_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg458_out;
SharedReg312_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg312_out;
SharedReg584_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg584_out;
SharedReg973_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg973_out;
SharedReg146_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg146_out;
SharedReg206_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg206_out;
SharedReg558_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg558_out;
SharedReg520_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg520_out;
SharedReg18_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg18_out;
SharedReg953_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg953_out;
SharedReg973_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg973_out;
SharedReg637_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg637_out;
   MUX_Subtract3_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg458_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg312_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg973_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg637_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg584_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg973_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg146_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg206_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg558_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg520_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg18_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg953_out_to_MUX_Subtract3_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract3_4_impl_1_out);

   Delay1No271_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_4_impl_1_out,
                 Y => Delay1No271_out);

Delay1No272_out_to_Subtract3_5_impl_parent_implementedSystem_port_0_cast <= Delay1No272_out;
Delay1No273_out_to_Subtract3_5_impl_parent_implementedSystem_port_1_cast <= Delay1No273_out;
   Subtract3_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract3_5_impl_out,
                 X => Delay1No272_out_to_Subtract3_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No273_out_to_Subtract3_5_impl_parent_implementedSystem_port_1_cast);

SharedReg904_out_to_MUX_Subtract3_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg904_out;
SharedReg903_out_to_MUX_Subtract3_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg903_out;
SharedReg903_out_to_MUX_Subtract3_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg903_out;
SharedReg1030_out_to_MUX_Subtract3_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1030_out;
SharedReg660_out_to_MUX_Subtract3_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg660_out;
SharedReg904_out_to_MUX_Subtract3_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg904_out;
SharedReg712_out_to_MUX_Subtract3_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg712_out;
SharedReg119_out_to_MUX_Subtract3_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg119_out;
SharedReg495_out_to_MUX_Subtract3_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg495_out;
Delay4No215_out_to_MUX_Subtract3_5_impl_0_parent_implementedSystem_port_10_cast <= Delay4No215_out;
SharedReg3_out_to_MUX_Subtract3_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg3_out;
SharedReg955_out_to_MUX_Subtract3_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg955_out;
   MUX_Subtract3_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg904_out_to_MUX_Subtract3_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg903_out_to_MUX_Subtract3_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg3_out_to_MUX_Subtract3_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg955_out_to_MUX_Subtract3_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg903_out_to_MUX_Subtract3_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1030_out_to_MUX_Subtract3_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg660_out_to_MUX_Subtract3_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg904_out_to_MUX_Subtract3_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg712_out_to_MUX_Subtract3_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg119_out_to_MUX_Subtract3_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg495_out_to_MUX_Subtract3_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay4No215_out_to_MUX_Subtract3_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract3_5_impl_0_out);

   Delay1No272_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_5_impl_0_out,
                 Y => Delay1No272_out);

SharedReg976_out_to_MUX_Subtract3_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg976_out;
SharedReg975_out_to_MUX_Subtract3_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg975_out;
SharedReg975_out_to_MUX_Subtract3_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg975_out;
SharedReg472_out_to_MUX_Subtract3_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg472_out;
SharedReg841_out_to_MUX_Subtract3_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg841_out;
SharedReg976_out_to_MUX_Subtract3_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg976_out;
SharedReg713_out_to_MUX_Subtract3_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg713_out;
SharedReg286_out_to_MUX_Subtract3_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg286_out;
SharedReg560_out_to_MUX_Subtract3_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg560_out;
SharedReg524_out_to_MUX_Subtract3_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg524_out;
SharedReg19_out_to_MUX_Subtract3_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg19_out;
SharedReg956_out_to_MUX_Subtract3_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg956_out;
   MUX_Subtract3_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg976_out_to_MUX_Subtract3_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg975_out_to_MUX_Subtract3_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg19_out_to_MUX_Subtract3_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg956_out_to_MUX_Subtract3_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg975_out_to_MUX_Subtract3_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg472_out_to_MUX_Subtract3_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg841_out_to_MUX_Subtract3_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg976_out_to_MUX_Subtract3_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg713_out_to_MUX_Subtract3_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg286_out_to_MUX_Subtract3_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg560_out_to_MUX_Subtract3_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg524_out_to_MUX_Subtract3_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract3_5_impl_1_out);

   Delay1No273_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_5_impl_1_out,
                 Y => Delay1No273_out);

Delay1No274_out_to_Subtract3_6_impl_parent_implementedSystem_port_0_cast <= Delay1No274_out;
Delay1No275_out_to_Subtract3_6_impl_parent_implementedSystem_port_1_cast <= Delay1No275_out;
   Subtract3_6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract3_6_impl_out,
                 X => Delay1No274_out_to_Subtract3_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No275_out_to_Subtract3_6_impl_parent_implementedSystem_port_1_cast);

SharedReg664_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg664_out;
SharedReg414_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg414_out;
SharedReg663_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg663_out;
SharedReg547_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg547_out;
SharedReg547_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg547_out;
SharedReg547_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg547_out;
SharedReg498_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg498_out;
SharedReg473_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg473_out;
SharedReg642_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg642_out;
SharedReg498_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg498_out;
SharedReg547_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg547_out;
SharedReg1_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1_out;
   MUX_Subtract3_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg664_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg414_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg547_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg663_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg547_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg547_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg547_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg498_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg473_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg642_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg498_out_to_MUX_Subtract3_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract3_6_impl_0_out);

   Delay1No274_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_6_impl_0_out,
                 Y => Delay1No274_out);

SharedReg846_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg846_out;
SharedReg526_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg526_out;
SharedReg845_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg845_out;
SharedReg642_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg642_out;
SharedReg642_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg642_out;
SharedReg642_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg642_out;
SharedReg562_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg562_out;
SharedReg700_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg700_out;
SharedReg818_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg818_out;
SharedReg562_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg562_out;
SharedReg642_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg642_out;
SharedReg17_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg17_out;
   MUX_Subtract3_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg846_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg526_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg642_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg17_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg845_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg642_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg642_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg642_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg562_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg700_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg818_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg562_out_to_MUX_Subtract3_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract3_6_impl_1_out);

   Delay1No275_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_6_impl_1_out,
                 Y => Delay1No275_out);

Delay1No276_out_to_Product6_0_impl_parent_implementedSystem_port_0_cast <= Delay1No276_out;
Delay1No277_out_to_Product6_0_impl_parent_implementedSystem_port_1_cast <= Delay1No277_out;
   Product6_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product6_0_impl_out,
                 X => Delay1No276_out_to_Product6_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No277_out_to_Product6_0_impl_parent_implementedSystem_port_1_cast);

SharedReg1120_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1120_out;
SharedReg1121_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1121_out;
SharedReg1140_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1140_out;
SharedReg1124_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1124_out;
SharedReg1110_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1110_out;
SharedReg1126_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1126_out;
SharedReg775_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg775_out;
SharedReg1128_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1128_out;
SharedReg1138_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1138_out;
SharedReg1106_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1106_out;
SharedReg1119_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1125_out;
   MUX_Product6_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1120_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1121_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1119_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1125_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1140_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1124_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1110_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1126_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg775_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1128_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1138_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1106_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product6_0_impl_0_out);

   Delay1No276_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_0_impl_0_out,
                 Y => Delay1No276_out);

SharedReg65_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg65_out;
SharedReg33_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg33_out;
SharedReg564_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg564_out;
SharedReg95_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg95_out;
SharedReg68_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg68_out;
SharedReg205_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg205_out;
SharedReg1156_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1156_out;
SharedReg982_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg982_out;
SharedReg1005_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1005_out;
SharedReg97_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg97_out;
SharedReg95_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg95_out;
SharedReg35_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg35_out;
   MUX_Product6_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg65_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg33_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg95_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg35_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg564_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg95_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg68_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg205_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1156_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg982_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1005_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg97_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product6_0_impl_1_out);

   Delay1No277_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_0_impl_1_out,
                 Y => Delay1No277_out);

Delay1No278_out_to_Product6_1_impl_parent_implementedSystem_port_0_cast <= Delay1No278_out;
Delay1No279_out_to_Product6_1_impl_parent_implementedSystem_port_1_cast <= Delay1No279_out;
   Product6_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product6_1_impl_out,
                 X => Delay1No278_out_to_Product6_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No279_out_to_Product6_1_impl_parent_implementedSystem_port_1_cast);

SharedReg1119_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1125_out;
SharedReg1120_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1120_out;
SharedReg1121_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1121_out;
SharedReg1140_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1140_out;
SharedReg1124_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1124_out;
SharedReg1110_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1110_out;
SharedReg1126_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1126_out;
SharedReg746_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg746_out;
SharedReg1128_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1128_out;
SharedReg1138_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1138_out;
SharedReg1106_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1106_out;
   MUX_Product6_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1119_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1125_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1138_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1106_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1120_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1121_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1140_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1124_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1110_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1126_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg746_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1128_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product6_1_impl_0_out);

   Delay1No278_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_1_impl_0_out,
                 Y => Delay1No278_out);

SharedReg69_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg69_out;
SharedReg161_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg161_out;
SharedReg38_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg38_out;
SharedReg159_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg159_out;
SharedReg438_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg438_out;
SharedReg69_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg69_out;
SharedReg40_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg40_out;
SharedReg133_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg133_out;
SharedReg1156_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1156_out;
SharedReg985_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg985_out;
SharedReg1008_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1008_out;
SharedReg102_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg102_out;
   MUX_Product6_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg69_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg161_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1008_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg102_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg38_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg159_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg438_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg69_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg40_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg133_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1156_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg985_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product6_1_impl_1_out);

   Delay1No279_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_1_impl_1_out,
                 Y => Delay1No279_out);

Delay1No280_out_to_Product6_2_impl_parent_implementedSystem_port_0_cast <= Delay1No280_out;
Delay1No281_out_to_Product6_2_impl_parent_implementedSystem_port_1_cast <= Delay1No281_out;
   Product6_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product6_2_impl_out,
                 X => Delay1No280_out_to_Product6_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No281_out_to_Product6_2_impl_parent_implementedSystem_port_1_cast);

SharedReg1138_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1138_out;
SharedReg1106_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1106_out;
SharedReg1119_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1125_out;
SharedReg1120_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1120_out;
SharedReg1121_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1121_out;
SharedReg1140_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1140_out;
SharedReg1124_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1124_out;
SharedReg1110_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1110_out;
SharedReg1126_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1126_out;
SharedReg753_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg753_out;
SharedReg1128_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1128_out;
   MUX_Product6_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1138_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1106_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg753_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1128_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1119_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1125_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1120_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1121_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1140_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1124_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1110_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1126_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product6_2_impl_0_out);

   Delay1No280_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_2_impl_0_out,
                 Y => Delay1No280_out);

SharedReg987_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg987_out;
SharedReg107_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg107_out;
SharedReg73_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg73_out;
SharedReg166_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg166_out;
SharedReg41_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg41_out;
SharedReg165_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg165_out;
SharedReg445_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg445_out;
SharedReg105_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg105_out;
SharedReg43_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg43_out;
SharedReg138_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg138_out;
SharedReg1156_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1156_out;
SharedReg859_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg859_out;
   MUX_Product6_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg987_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg107_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1156_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg859_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg73_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg166_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg41_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg165_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg445_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg105_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg43_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg138_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product6_2_impl_1_out);

   Delay1No281_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_2_impl_1_out,
                 Y => Delay1No281_out);

Delay1No282_out_to_Product6_3_impl_parent_implementedSystem_port_0_cast <= Delay1No282_out;
Delay1No283_out_to_Product6_3_impl_parent_implementedSystem_port_1_cast <= Delay1No283_out;
   Product6_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product6_3_impl_out,
                 X => Delay1No282_out_to_Product6_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No283_out_to_Product6_3_impl_parent_implementedSystem_port_1_cast);

SharedReg1128_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1128_out;
SharedReg1138_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1138_out;
SharedReg1106_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1106_out;
SharedReg1119_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1125_out;
SharedReg1120_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1120_out;
SharedReg1121_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1121_out;
SharedReg1140_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1140_out;
SharedReg1124_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1124_out;
SharedReg1110_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1110_out;
SharedReg1126_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1126_out;
SharedReg705_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg705_out;
   MUX_Product6_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1128_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1138_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1126_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg705_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1106_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1119_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1125_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1120_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1121_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1140_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1124_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1110_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product6_3_impl_0_out);

   Delay1No282_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_3_impl_0_out,
                 Y => Delay1No282_out);

SharedReg991_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg991_out;
SharedReg991_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg991_out;
SharedReg79_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg79_out;
SharedReg44_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg44_out;
SharedReg200_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg200_out;
SharedReg198_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg198_out;
SharedReg171_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg171_out;
SharedReg451_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg451_out;
SharedReg110_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg110_out;
SharedReg47_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg47_out;
SharedReg113_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg113_out;
SharedReg1156_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1156_out;
   MUX_Product6_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg991_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg991_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg113_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1156_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg79_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg44_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg200_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg198_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg171_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg451_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg110_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg47_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product6_3_impl_1_out);

   Delay1No283_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_3_impl_1_out,
                 Y => Delay1No283_out);

Delay1No284_out_to_Product6_4_impl_parent_implementedSystem_port_0_cast <= Delay1No284_out;
Delay1No285_out_to_Product6_4_impl_parent_implementedSystem_port_1_cast <= Delay1No285_out;
   Product6_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product6_4_impl_out,
                 X => Delay1No284_out_to_Product6_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No285_out_to_Product6_4_impl_parent_implementedSystem_port_1_cast);

SharedReg1126_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1126_out;
SharedReg712_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg712_out;
SharedReg1128_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1128_out;
SharedReg1138_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1138_out;
SharedReg1106_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1106_out;
SharedReg1119_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1125_out;
SharedReg1120_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1120_out;
SharedReg1121_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1121_out;
SharedReg1140_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1140_out;
SharedReg1124_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1124_out;
SharedReg1110_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1110_out;
   MUX_Product6_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1126_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg712_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1124_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1110_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1128_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1138_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1106_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1119_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1125_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1120_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1121_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1140_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product6_4_impl_0_out);

   Delay1No284_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_4_impl_0_out,
                 Y => Delay1No284_out);

SharedReg117_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg117_out;
SharedReg1156_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1156_out;
SharedReg866_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg866_out;
SharedReg866_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg866_out;
SharedReg83_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg83_out;
SharedReg48_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg48_out;
SharedReg193_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg193_out;
SharedReg48_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg48_out;
SharedReg176_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg176_out;
SharedReg458_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg458_out;
SharedReg114_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg114_out;
SharedReg84_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg84_out;
   MUX_Product6_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg117_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1156_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg114_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg84_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg866_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg866_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg83_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg48_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg193_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg48_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg176_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg458_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product6_4_impl_1_out);

   Delay1No285_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_4_impl_1_out,
                 Y => Delay1No285_out);

Delay1No286_out_to_Product6_5_impl_parent_implementedSystem_port_0_cast <= Delay1No286_out;
Delay1No287_out_to_Product6_5_impl_parent_implementedSystem_port_1_cast <= Delay1No287_out;
   Product6_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product6_5_impl_out,
                 X => Delay1No286_out_to_Product6_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No287_out_to_Product6_5_impl_parent_implementedSystem_port_1_cast);

SharedReg1124_out_to_MUX_Product6_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1124_out;
SharedReg1110_out_to_MUX_Product6_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1110_out;
SharedReg1126_out_to_MUX_Product6_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1126_out;
SharedReg770_out_to_MUX_Product6_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg770_out;
SharedReg1128_out_to_MUX_Product6_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1128_out;
SharedReg1138_out_to_MUX_Product6_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1138_out;
SharedReg1106_out_to_MUX_Product6_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1106_out;
SharedReg1119_out_to_MUX_Product6_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product6_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1125_out;
SharedReg1120_out_to_MUX_Product6_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1120_out;
SharedReg1121_out_to_MUX_Product6_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1121_out;
SharedReg1140_out_to_MUX_Product6_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1140_out;
   MUX_Product6_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1124_out_to_MUX_Product6_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1110_out_to_MUX_Product6_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1121_out_to_MUX_Product6_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1140_out_to_MUX_Product6_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1126_out_to_MUX_Product6_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg770_out_to_MUX_Product6_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1128_out_to_MUX_Product6_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1138_out_to_MUX_Product6_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1106_out_to_MUX_Product6_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1119_out_to_MUX_Product6_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1125_out_to_MUX_Product6_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1120_out_to_MUX_Product6_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product6_5_impl_0_out);

   Delay1No286_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_5_impl_0_out,
                 Y => Delay1No286_out);

SharedReg150_out_to_MUX_Product6_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg150_out;
SharedReg121_out_to_MUX_Product6_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg121_out;
SharedReg186_out_to_MUX_Product6_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg186_out;
SharedReg1156_out_to_MUX_Product6_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1156_out;
SharedReg695_out_to_MUX_Product6_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg695_out;
SharedReg869_out_to_MUX_Product6_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg869_out;
SharedReg120_out_to_MUX_Product6_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg120_out;
SharedReg118_out_to_MUX_Product6_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg118_out;
SharedReg281_out_to_MUX_Product6_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg281_out;
SharedReg118_out_to_MUX_Product6_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg118_out;
SharedReg87_out_to_MUX_Product6_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg87_out;
SharedReg589_out_to_MUX_Product6_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg589_out;
   MUX_Product6_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg150_out_to_MUX_Product6_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg121_out_to_MUX_Product6_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg87_out_to_MUX_Product6_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg589_out_to_MUX_Product6_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg186_out_to_MUX_Product6_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1156_out_to_MUX_Product6_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg695_out_to_MUX_Product6_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg869_out_to_MUX_Product6_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg120_out_to_MUX_Product6_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg118_out_to_MUX_Product6_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg281_out_to_MUX_Product6_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg118_out_to_MUX_Product6_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product6_5_impl_1_out);

   Delay1No287_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_5_impl_1_out,
                 Y => Delay1No287_out);

Delay1No288_out_to_Product6_6_impl_parent_implementedSystem_port_0_cast <= Delay1No288_out;
Delay1No289_out_to_Product6_6_impl_parent_implementedSystem_port_1_cast <= Delay1No289_out;
   Product6_6_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product6_6_impl_out,
                 X => Delay1No288_out_to_Product6_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No289_out_to_Product6_6_impl_parent_implementedSystem_port_1_cast);

SharedReg1140_out_to_MUX_Product6_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1140_out;
SharedReg1124_out_to_MUX_Product6_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1124_out;
SharedReg1110_out_to_MUX_Product6_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1110_out;
SharedReg1126_out_to_MUX_Product6_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1126_out;
SharedReg1101_out_to_MUX_Product6_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1101_out;
SharedReg1128_out_to_MUX_Product6_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1128_out;
SharedReg1138_out_to_MUX_Product6_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1138_out;
SharedReg1106_out_to_MUX_Product6_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1106_out;
SharedReg1119_out_to_MUX_Product6_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product6_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1125_out;
SharedReg1120_out_to_MUX_Product6_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1120_out;
SharedReg1121_out_to_MUX_Product6_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1121_out;
   MUX_Product6_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1140_out_to_MUX_Product6_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1124_out_to_MUX_Product6_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1120_out_to_MUX_Product6_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1121_out_to_MUX_Product6_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1110_out_to_MUX_Product6_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1126_out_to_MUX_Product6_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1101_out_to_MUX_Product6_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1128_out_to_MUX_Product6_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1138_out_to_MUX_Product6_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1106_out_to_MUX_Product6_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1119_out_to_MUX_Product6_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1125_out_to_MUX_Product6_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product6_6_impl_0_out);

   Delay1No288_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_6_impl_0_out,
                 Y => Delay1No288_out);

SharedReg595_out_to_MUX_Product6_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg595_out;
SharedReg153_out_to_MUX_Product6_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg153_out;
SharedReg125_out_to_MUX_Product6_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg125_out;
SharedReg190_out_to_MUX_Product6_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg190_out;
SharedReg1156_out_to_MUX_Product6_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1156_out;
SharedReg1002_out_to_MUX_Product6_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1002_out;
SharedReg1002_out_to_MUX_Product6_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1002_out;
SharedReg93_out_to_MUX_Product6_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg93_out;
SharedReg123_out_to_MUX_Product6_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg123_out;
SharedReg63_out_to_MUX_Product6_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg63_out;
SharedReg91_out_to_MUX_Product6_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg91_out;
SharedReg61_out_to_MUX_Product6_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg61_out;
   MUX_Product6_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg595_out_to_MUX_Product6_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg153_out_to_MUX_Product6_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg91_out_to_MUX_Product6_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg61_out_to_MUX_Product6_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg125_out_to_MUX_Product6_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg190_out_to_MUX_Product6_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1156_out_to_MUX_Product6_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1002_out_to_MUX_Product6_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1002_out_to_MUX_Product6_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg93_out_to_MUX_Product6_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg123_out_to_MUX_Product6_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg63_out_to_MUX_Product6_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product6_6_impl_1_out);

   Delay1No289_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_6_impl_1_out,
                 Y => Delay1No289_out);

Delay1No290_out_to_Product23_0_impl_parent_implementedSystem_port_0_cast <= Delay1No290_out;
Delay1No291_out_to_Product23_0_impl_parent_implementedSystem_port_1_cast <= Delay1No291_out;
   Product23_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product23_0_impl_out,
                 X => Delay1No290_out_to_Product23_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No291_out_to_Product23_0_impl_parent_implementedSystem_port_1_cast);

SharedReg95_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg95_out;
SharedReg127_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg127_out;
SharedReg666_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg666_out;
SharedReg127_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg127_out;
SharedReg1110_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1110_out;
SharedReg36_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg36_out;
SharedReg1103_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1103_out;
SharedReg1130_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1130_out;
SharedReg1038_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1038_out;
SharedReg1118_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1118_out;
SharedReg127_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg127_out;
SharedReg68_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg68_out;
   MUX_Product23_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg95_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg127_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg127_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg68_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg666_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg127_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1110_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg36_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1103_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1130_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1038_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1118_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product23_0_impl_0_out);

   Delay1No290_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_0_impl_0_out,
                 Y => Delay1No290_out);

SharedReg1120_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1120_out;
SharedReg1121_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1121_out;
SharedReg1140_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1140_out;
SharedReg1124_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1124_out;
SharedReg98_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg98_out;
SharedReg1126_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1126_out;
SharedReg202_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg202_out;
SharedReg982_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg982_out;
SharedReg1138_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1138_out;
SharedReg97_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg97_out;
SharedReg1119_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1125_out;
   MUX_Product23_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1120_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1121_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1119_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1125_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1140_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1124_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg98_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1126_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg202_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg982_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1138_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg97_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product23_0_impl_1_out);

   Delay1No291_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_0_impl_1_out,
                 Y => Delay1No291_out);

Delay1No292_out_to_Product23_1_impl_parent_implementedSystem_port_0_cast <= Delay1No292_out;
Delay1No293_out_to_Product23_1_impl_parent_implementedSystem_port_1_cast <= Delay1No293_out;
   Product23_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product23_1_impl_out,
                 X => Delay1No292_out_to_Product23_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No293_out_to_Product23_1_impl_parent_implementedSystem_port_1_cast);

SharedReg100_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg100_out;
SharedReg40_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg40_out;
SharedReg69_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg69_out;
SharedReg100_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg100_out;
SharedReg570_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg570_out;
SharedReg100_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg100_out;
SharedReg1110_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1110_out;
SharedReg162_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg162_out;
SharedReg1103_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1103_out;
SharedReg1130_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1130_out;
SharedReg1043_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1043_out;
SharedReg1118_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1118_out;
   MUX_Product23_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg100_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg40_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1043_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1118_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg69_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg100_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg570_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg100_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1110_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg162_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1103_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1130_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product23_1_impl_0_out);

   Delay1No292_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_1_impl_0_out,
                 Y => Delay1No292_out);

SharedReg1119_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1125_out;
SharedReg1120_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1120_out;
SharedReg1121_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1121_out;
SharedReg1140_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1140_out;
SharedReg1124_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1124_out;
SharedReg72_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg72_out;
SharedReg1126_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1126_out;
SharedReg234_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg234_out;
SharedReg985_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg985_out;
SharedReg1138_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1138_out;
SharedReg102_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg102_out;
   MUX_Product23_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1119_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1125_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1138_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg102_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1120_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1121_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1140_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1124_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg72_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1126_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg234_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg985_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product23_1_impl_1_out);

   Delay1No293_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_1_impl_1_out,
                 Y => Delay1No293_out);

Delay1No294_out_to_Product23_2_impl_parent_implementedSystem_port_0_cast <= Delay1No294_out;
Delay1No295_out_to_Product23_2_impl_parent_implementedSystem_port_1_cast <= Delay1No295_out;
   Product23_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product23_2_impl_out,
                 X => Delay1No294_out_to_Product23_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No295_out_to_Product23_2_impl_parent_implementedSystem_port_1_cast);

SharedReg1013_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1013_out;
SharedReg1118_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1118_out;
SharedReg105_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg105_out;
SharedReg43_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg43_out;
SharedReg73_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg73_out;
SharedReg105_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg105_out;
SharedReg576_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg576_out;
SharedReg134_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg134_out;
SharedReg1110_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1110_out;
SharedReg167_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg167_out;
SharedReg1103_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1103_out;
SharedReg1130_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1130_out;
   MUX_Product23_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1013_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1118_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1103_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1130_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg105_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg43_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg73_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg105_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg576_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg134_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1110_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg167_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product23_2_impl_0_out);

   Delay1No294_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_2_impl_0_out,
                 Y => Delay1No294_out);

SharedReg1138_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1138_out;
SharedReg107_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg107_out;
SharedReg1119_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1125_out;
SharedReg1120_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1120_out;
SharedReg1121_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1121_out;
SharedReg1140_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1140_out;
SharedReg1124_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1124_out;
SharedReg76_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg76_out;
SharedReg1126_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1126_out;
SharedReg239_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg239_out;
SharedReg859_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg859_out;
   MUX_Product23_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1138_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg107_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg239_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg859_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1119_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1125_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1120_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1121_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1140_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1124_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg76_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1126_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product23_2_impl_1_out);

   Delay1No295_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_2_impl_1_out,
                 Y => Delay1No295_out);

Delay1No296_out_to_Product23_3_impl_parent_implementedSystem_port_0_cast <= Delay1No296_out;
Delay1No297_out_to_Product23_3_impl_parent_implementedSystem_port_1_cast <= Delay1No297_out;
   Product23_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product23_3_impl_out,
                 X => Delay1No296_out_to_Product23_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No297_out_to_Product23_3_impl_parent_implementedSystem_port_1_cast);

SharedReg1130_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1130_out;
SharedReg1018_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1018_out;
SharedReg1118_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1118_out;
SharedReg77_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg77_out;
SharedReg47_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg47_out;
SharedReg44_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg44_out;
SharedReg110_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg110_out;
SharedReg580_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg580_out;
SharedReg139_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg139_out;
SharedReg1110_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1110_out;
SharedReg172_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg172_out;
SharedReg1103_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1103_out;
   MUX_Product23_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1130_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1018_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg172_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1103_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1118_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg77_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg47_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg44_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg110_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg580_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg139_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1110_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product23_3_impl_0_out);

   Delay1No296_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_3_impl_0_out,
                 Y => Delay1No296_out);

SharedReg991_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg991_out;
SharedReg1138_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1138_out;
SharedReg79_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg79_out;
SharedReg1119_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1125_out;
SharedReg1120_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1120_out;
SharedReg1121_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1121_out;
SharedReg1140_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1140_out;
SharedReg1124_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1124_out;
SharedReg80_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg80_out;
SharedReg1126_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1126_out;
SharedReg244_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg244_out;
   MUX_Product23_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg991_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1138_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1126_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg244_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg79_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1119_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1125_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1120_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1121_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1140_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1124_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg80_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product23_3_impl_1_out);

   Delay1No297_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_3_impl_1_out,
                 Y => Delay1No297_out);

Delay1No298_out_to_Product23_4_impl_parent_implementedSystem_port_0_cast <= Delay1No298_out;
Delay1No299_out_to_Product23_4_impl_parent_implementedSystem_port_1_cast <= Delay1No299_out;
   Product23_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product23_4_impl_out,
                 X => Delay1No298_out_to_Product23_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No299_out_to_Product23_4_impl_parent_implementedSystem_port_1_cast);

SharedReg179_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg179_out;
SharedReg1103_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1103_out;
SharedReg1130_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1130_out;
SharedReg994_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg994_out;
SharedReg1118_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1118_out;
SharedReg81_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg81_out;
SharedReg178_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg178_out;
SharedReg81_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg81_out;
SharedReg145_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg145_out;
SharedReg584_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg584_out;
SharedReg145_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg145_out;
SharedReg1110_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1110_out;
   MUX_Product23_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg179_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1103_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg145_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1110_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1130_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg994_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1118_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg81_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg178_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg81_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg145_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg584_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product23_4_impl_0_out);

   Delay1No298_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_4_impl_0_out,
                 Y => Delay1No298_out);

SharedReg1126_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1126_out;
SharedReg206_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg206_out;
SharedReg866_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg866_out;
SharedReg1138_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1138_out;
SharedReg83_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg83_out;
SharedReg1119_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1125_out;
SharedReg1120_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1120_out;
SharedReg1121_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1121_out;
SharedReg1140_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1140_out;
SharedReg1124_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1124_out;
SharedReg116_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg116_out;
   MUX_Product23_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1126_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg206_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1124_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg116_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg866_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1138_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg83_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1119_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1125_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1120_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1121_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1140_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product23_4_impl_1_out);

   Delay1No299_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_4_impl_1_out,
                 Y => Delay1No299_out);

Delay1No300_out_to_Product23_5_impl_parent_implementedSystem_port_0_cast <= Delay1No300_out;
Delay1No301_out_to_Product23_5_impl_parent_implementedSystem_port_1_cast <= Delay1No301_out;
   Product23_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product23_5_impl_out,
                 X => Delay1No300_out_to_Product23_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No301_out_to_Product23_5_impl_parent_implementedSystem_port_1_cast);

SharedReg182_out_to_MUX_Product23_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg182_out;
SharedReg1110_out_to_MUX_Product23_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1110_out;
SharedReg90_out_to_MUX_Product23_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg90_out;
SharedReg1103_out_to_MUX_Product23_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1103_out;
SharedReg1130_out_to_MUX_Product23_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1130_out;
SharedReg998_out_to_MUX_Product23_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg998_out;
SharedReg1118_out_to_MUX_Product23_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1118_out;
SharedReg150_out_to_MUX_Product23_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg150_out;
SharedReg55_out_to_MUX_Product23_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg55_out;
SharedReg150_out_to_MUX_Product23_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg150_out;
SharedReg182_out_to_MUX_Product23_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg182_out;
SharedReg694_out_to_MUX_Product23_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg694_out;
   MUX_Product23_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg182_out_to_MUX_Product23_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1110_out_to_MUX_Product23_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg182_out_to_MUX_Product23_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg694_out_to_MUX_Product23_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg90_out_to_MUX_Product23_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1103_out_to_MUX_Product23_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1130_out_to_MUX_Product23_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg998_out_to_MUX_Product23_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1118_out_to_MUX_Product23_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg150_out_to_MUX_Product23_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg55_out_to_MUX_Product23_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg150_out_to_MUX_Product23_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product23_5_impl_0_out);

   Delay1No300_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_5_impl_0_out,
                 Y => Delay1No300_out);

SharedReg1124_out_to_MUX_Product23_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1124_out;
SharedReg152_out_to_MUX_Product23_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg152_out;
SharedReg1126_out_to_MUX_Product23_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1126_out;
SharedReg182_out_to_MUX_Product23_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg182_out;
SharedReg695_out_to_MUX_Product23_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg695_out;
SharedReg1138_out_to_MUX_Product23_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1138_out;
SharedReg120_out_to_MUX_Product23_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg120_out;
SharedReg1119_out_to_MUX_Product23_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product23_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1125_out;
SharedReg1120_out_to_MUX_Product23_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1120_out;
SharedReg1121_out_to_MUX_Product23_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1121_out;
SharedReg1140_out_to_MUX_Product23_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1140_out;
   MUX_Product23_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1124_out_to_MUX_Product23_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg152_out_to_MUX_Product23_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1121_out_to_MUX_Product23_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1140_out_to_MUX_Product23_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1126_out_to_MUX_Product23_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg182_out_to_MUX_Product23_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg695_out_to_MUX_Product23_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1138_out_to_MUX_Product23_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg120_out_to_MUX_Product23_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1119_out_to_MUX_Product23_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1125_out_to_MUX_Product23_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1120_out_to_MUX_Product23_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product23_5_impl_1_out);

   Delay1No301_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_5_impl_1_out,
                 Y => Delay1No301_out);

Delay1No302_out_to_Product23_6_impl_parent_implementedSystem_port_0_cast <= Delay1No302_out;
Delay1No303_out_to_Product23_6_impl_parent_implementedSystem_port_1_cast <= Delay1No303_out;
   Product23_6_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product23_6_impl_out,
                 X => Delay1No302_out_to_Product23_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No303_out_to_Product23_6_impl_parent_implementedSystem_port_1_cast);

SharedReg699_out_to_MUX_Product23_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg699_out;
SharedReg187_out_to_MUX_Product23_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg187_out;
SharedReg1110_out_to_MUX_Product23_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1110_out;
SharedReg64_out_to_MUX_Product23_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg64_out;
SharedReg1103_out_to_MUX_Product23_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1103_out;
SharedReg1130_out_to_MUX_Product23_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1130_out;
SharedReg1034_out_to_MUX_Product23_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1034_out;
SharedReg1118_out_to_MUX_Product23_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1118_out;
SharedReg153_out_to_MUX_Product23_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg153_out;
SharedReg94_out_to_MUX_Product23_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg94_out;
SharedReg123_out_to_MUX_Product23_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg123_out;
SharedReg187_out_to_MUX_Product23_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg187_out;
   MUX_Product23_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg699_out_to_MUX_Product23_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg187_out_to_MUX_Product23_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg123_out_to_MUX_Product23_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg187_out_to_MUX_Product23_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1110_out_to_MUX_Product23_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg64_out_to_MUX_Product23_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1103_out_to_MUX_Product23_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1130_out_to_MUX_Product23_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1034_out_to_MUX_Product23_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1118_out_to_MUX_Product23_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg153_out_to_MUX_Product23_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg94_out_to_MUX_Product23_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product23_6_impl_0_out);

   Delay1No302_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_6_impl_0_out,
                 Y => Delay1No302_out);

SharedReg1140_out_to_MUX_Product23_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1140_out;
SharedReg1124_out_to_MUX_Product23_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1124_out;
SharedReg156_out_to_MUX_Product23_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg156_out;
SharedReg1126_out_to_MUX_Product23_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1126_out;
SharedReg187_out_to_MUX_Product23_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg187_out;
SharedReg1002_out_to_MUX_Product23_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1002_out;
SharedReg1138_out_to_MUX_Product23_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1138_out;
SharedReg93_out_to_MUX_Product23_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg93_out;
SharedReg1119_out_to_MUX_Product23_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product23_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1125_out;
SharedReg1120_out_to_MUX_Product23_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1120_out;
SharedReg1121_out_to_MUX_Product23_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1121_out;
   MUX_Product23_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1140_out_to_MUX_Product23_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1124_out_to_MUX_Product23_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1120_out_to_MUX_Product23_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1121_out_to_MUX_Product23_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg156_out_to_MUX_Product23_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1126_out_to_MUX_Product23_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg187_out_to_MUX_Product23_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1002_out_to_MUX_Product23_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1138_out_to_MUX_Product23_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg93_out_to_MUX_Product23_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1119_out_to_MUX_Product23_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1125_out_to_MUX_Product23_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product23_6_impl_1_out);

   Delay1No303_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_6_impl_1_out,
                 Y => Delay1No303_out);

Delay1No304_out_to_Product33_0_impl_parent_implementedSystem_port_0_cast <= Delay1No304_out;
Delay1No305_out_to_Product33_0_impl_parent_implementedSystem_port_1_cast <= Delay1No305_out;
   Product33_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product33_0_impl_out,
                 X => Delay1No304_out_to_Product33_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No305_out_to_Product33_0_impl_parent_implementedSystem_port_1_cast);

SharedReg1129_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1129_out;
SharedReg1109_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1109_out;
SharedReg1111_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1111_out;
SharedReg1137_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1137_out;
SharedReg1135_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1135_out;
SharedReg1114_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1114_out;
SharedReg1103_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1103_out;
SharedReg1005_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1005_out;
SharedReg1142_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1142_out;
SharedReg1106_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1106_out;
SharedReg1107_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1113_out;
   MUX_Product33_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1129_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1109_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1107_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1113_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1111_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1137_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1135_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1114_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1103_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1005_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1142_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1106_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product33_0_impl_0_out);

   Delay1No304_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_0_impl_0_out,
                 Y => Delay1No304_out);

SharedReg981_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg981_out;
SharedReg1094_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1094_out;
SharedReg32_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg32_out;
SharedReg849_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg849_out;
SharedReg851_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg851_out;
SharedReg1099_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1099_out;
SharedReg249_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg249_out;
SharedReg1130_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1130_out;
SharedReg1072_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1072_out;
SharedReg329_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg329_out;
SharedReg981_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg981_out;
SharedReg1073_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1073_out;
   MUX_Product33_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg981_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1094_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg981_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1073_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg32_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg849_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg851_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1099_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg249_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1130_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1072_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg329_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product33_0_impl_1_out);

   Delay1No305_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_0_impl_1_out,
                 Y => Delay1No305_out);

Delay1No306_out_to_Product33_1_impl_parent_implementedSystem_port_0_cast <= Delay1No306_out;
Delay1No307_out_to_Product33_1_impl_parent_implementedSystem_port_1_cast <= Delay1No307_out;
   Product33_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product33_1_impl_out,
                 X => Delay1No306_out_to_Product33_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No307_out_to_Product33_1_impl_parent_implementedSystem_port_1_cast);

SharedReg1107_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1113_out;
SharedReg1129_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1129_out;
SharedReg1109_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1109_out;
SharedReg1111_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1111_out;
SharedReg1137_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1137_out;
SharedReg1135_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1135_out;
SharedReg1114_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1114_out;
SharedReg1103_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1103_out;
SharedReg1008_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1008_out;
SharedReg1142_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1142_out;
SharedReg1106_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1106_out;
   MUX_Product33_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1107_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1113_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1142_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1106_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1129_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1109_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1111_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1137_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1135_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1114_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1103_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1008_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product33_1_impl_0_out);

   Delay1No306_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_1_impl_0_out,
                 Y => Delay1No306_out);

SharedReg854_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg854_out;
SharedReg1045_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1045_out;
SharedReg854_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg854_out;
SharedReg1081_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1081_out;
SharedReg158_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg158_out;
SharedReg672_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg672_out;
SharedReg674_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg674_out;
SharedReg1086_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1086_out;
SharedReg254_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg254_out;
SharedReg1130_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1130_out;
SharedReg1083_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1083_out;
SharedReg374_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg374_out;
   MUX_Product33_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg854_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1045_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1083_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg374_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg854_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1081_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg158_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg672_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg674_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1086_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg254_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1130_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product33_1_impl_1_out);

   Delay1No307_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_1_impl_1_out,
                 Y => Delay1No307_out);

Delay1No308_out_to_Product33_2_impl_parent_implementedSystem_port_0_cast <= Delay1No308_out;
Delay1No309_out_to_Product33_2_impl_parent_implementedSystem_port_1_cast <= Delay1No309_out;
   Product33_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product33_2_impl_out,
                 X => Delay1No308_out_to_Product33_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No309_out_to_Product33_2_impl_parent_implementedSystem_port_1_cast);

SharedReg1142_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1142_out;
SharedReg1106_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1106_out;
SharedReg1107_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1113_out;
SharedReg1129_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1129_out;
SharedReg1109_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1109_out;
SharedReg1111_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1111_out;
SharedReg1137_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1137_out;
SharedReg1135_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1135_out;
SharedReg1114_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1114_out;
SharedReg1103_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1103_out;
SharedReg987_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg987_out;
   MUX_Product33_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1142_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1106_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1103_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg987_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1107_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1113_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1129_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1109_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1111_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1137_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1135_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1114_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product33_2_impl_0_out);

   Delay1No308_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_2_impl_0_out,
                 Y => Delay1No308_out);

SharedReg1049_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1049_out;
SharedReg345_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg345_out;
SharedReg678_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg678_out;
SharedReg1015_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1015_out;
SharedReg678_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg678_out;
SharedReg1047_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1047_out;
SharedReg41_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg41_out;
SharedReg678_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg678_out;
SharedReg578_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg578_out;
SharedReg1052_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1052_out;
SharedReg260_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg260_out;
SharedReg1130_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1130_out;
   MUX_Product33_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1049_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg345_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg260_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1130_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg678_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1015_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg678_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1047_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg41_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg678_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg578_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1052_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product33_2_impl_1_out);

   Delay1No309_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_2_impl_1_out,
                 Y => Delay1No309_out);

Delay1No310_out_to_Product33_3_impl_parent_implementedSystem_port_0_cast <= Delay1No310_out;
Delay1No311_out_to_Product33_3_impl_parent_implementedSystem_port_1_cast <= Delay1No311_out;
   Product33_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product33_3_impl_out,
                 X => Delay1No310_out_to_Product33_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No311_out_to_Product33_3_impl_parent_implementedSystem_port_1_cast);

SharedReg1018_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1018_out;
SharedReg1142_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1142_out;
SharedReg1106_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1106_out;
SharedReg1107_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1113_out;
SharedReg1129_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1129_out;
SharedReg1109_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1109_out;
SharedReg1111_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1111_out;
SharedReg1137_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1137_out;
SharedReg1135_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1135_out;
SharedReg1114_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1114_out;
SharedReg1103_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1103_out;
   MUX_Product33_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1018_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1142_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1114_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1103_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1106_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1107_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1113_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1129_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1109_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1111_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1137_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1135_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product33_3_impl_0_out);

   Delay1No310_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_3_impl_0_out,
                 Y => Delay1No310_out);

SharedReg1130_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1130_out;
SharedReg792_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg792_out;
SharedReg193_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg193_out;
SharedReg683_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg683_out;
SharedReg1056_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1056_out;
SharedReg683_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg683_out;
SharedReg790_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg790_out;
SharedReg198_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg198_out;
SharedReg861_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg861_out;
SharedReg685_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg685_out;
SharedReg1058_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1058_out;
SharedReg266_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg266_out;
   MUX_Product33_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1130_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg792_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1058_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg266_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg193_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg683_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1056_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg683_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg790_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg198_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg861_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg685_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product33_3_impl_1_out);

   Delay1No311_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_3_impl_1_out,
                 Y => Delay1No311_out);

Delay1No312_out_to_Product33_4_impl_parent_implementedSystem_port_0_cast <= Delay1No312_out;
Delay1No313_out_to_Product33_4_impl_parent_implementedSystem_port_1_cast <= Delay1No313_out;
   Product33_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product33_4_impl_out,
                 X => Delay1No312_out_to_Product33_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No313_out_to_Product33_4_impl_parent_implementedSystem_port_1_cast);

SharedReg1114_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1114_out;
SharedReg1103_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1103_out;
SharedReg994_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg994_out;
SharedReg1142_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1142_out;
SharedReg1106_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1106_out;
SharedReg1107_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1113_out;
SharedReg1129_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1129_out;
SharedReg1109_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1109_out;
SharedReg1111_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1111_out;
SharedReg1137_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1137_out;
SharedReg1135_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1135_out;
   MUX_Product33_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1114_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1103_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1137_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1135_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg994_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1142_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1106_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1107_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1113_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1129_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1109_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1111_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product33_4_impl_0_out);

   Delay1No312_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_4_impl_0_out,
                 Y => Delay1No312_out);

SharedReg1025_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1025_out;
SharedReg272_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg272_out;
SharedReg1130_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1130_out;
SharedReg797_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg797_out;
SharedReg281_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg281_out;
SharedReg584_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg584_out;
SharedReg995_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg995_out;
SharedReg689_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg689_out;
SharedReg764_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg764_out;
SharedReg48_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg48_out;
SharedReg689_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg689_out;
SharedReg691_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg691_out;
   MUX_Product33_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1025_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg272_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg689_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg691_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1130_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg797_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg281_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg584_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg995_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg689_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg764_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg48_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product33_4_impl_1_out);

   Delay1No313_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_4_impl_1_out,
                 Y => Delay1No313_out);

Delay1No314_out_to_Product33_5_impl_parent_implementedSystem_port_0_cast <= Delay1No314_out;
Delay1No315_out_to_Product33_5_impl_parent_implementedSystem_port_1_cast <= Delay1No315_out;
   Product33_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product33_5_impl_out,
                 X => Delay1No314_out_to_Product33_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No315_out_to_Product33_5_impl_parent_implementedSystem_port_1_cast);

SharedReg1137_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1137_out;
SharedReg1135_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1135_out;
SharedReg1114_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1114_out;
SharedReg1103_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1103_out;
SharedReg869_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg869_out;
SharedReg1142_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1142_out;
SharedReg1106_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1106_out;
SharedReg1107_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1113_out;
SharedReg1129_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1129_out;
SharedReg1109_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1109_out;
SharedReg1111_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1111_out;
   MUX_Product33_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1137_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1135_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1109_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1111_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1114_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1103_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg869_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1142_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1106_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1107_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1113_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1129_out_to_MUX_Product33_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product33_5_impl_0_out);

   Delay1No314_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_5_impl_0_out,
                 Y => Delay1No314_out);

SharedReg694_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg694_out;
SharedReg696_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg696_out;
SharedReg1063_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1063_out;
SharedReg212_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg212_out;
SharedReg1130_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1130_out;
SharedReg1030_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1030_out;
SharedReg293_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg293_out;
SharedReg694_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg694_out;
SharedReg1000_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1000_out;
SharedReg868_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg868_out;
SharedReg770_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg770_out;
SharedReg118_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg118_out;
   MUX_Product33_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg694_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg696_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg770_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg118_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1063_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg212_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1130_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1030_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg293_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg694_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1000_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg868_out_to_MUX_Product33_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product33_5_impl_1_out);

   Delay1No315_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_5_impl_1_out,
                 Y => Delay1No315_out);

Delay1No316_out_to_Product33_6_impl_parent_implementedSystem_port_0_cast <= Delay1No316_out;
Delay1No317_out_to_Product33_6_impl_parent_implementedSystem_port_1_cast <= Delay1No317_out;
   Product33_6_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product33_6_impl_out,
                 X => Delay1No316_out_to_Product33_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No317_out_to_Product33_6_impl_parent_implementedSystem_port_1_cast);

SharedReg1111_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1111_out;
SharedReg1137_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1137_out;
SharedReg1135_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1135_out;
SharedReg1114_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1114_out;
SharedReg1103_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1103_out;
SharedReg1034_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1034_out;
SharedReg1142_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1142_out;
SharedReg1106_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1106_out;
SharedReg1107_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1113_out;
SharedReg1129_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1129_out;
SharedReg1109_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1109_out;
   MUX_Product33_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1111_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1137_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1129_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1109_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1135_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1114_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1103_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1034_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1142_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1106_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1107_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1113_out_to_MUX_Product33_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product33_6_impl_0_out);

   Delay1No316_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_6_impl_0_out,
                 Y => Delay1No316_out);

SharedReg60_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg60_out;
SharedReg1001_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1001_out;
SharedReg1003_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1003_out;
SharedReg1093_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1093_out;
SharedReg218_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg218_out;
SharedReg1130_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1130_out;
SharedReg1077_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1077_out;
SharedReg358_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg358_out;
SharedReg1001_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1001_out;
SharedReg1078_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1078_out;
SharedReg1001_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1001_out;
SharedReg1101_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1101_out;
   MUX_Product33_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg60_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1001_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1001_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1101_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1003_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1093_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg218_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1130_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1077_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg358_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1001_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1078_out_to_MUX_Product33_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product33_6_impl_1_out);

   Delay1No317_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_6_impl_1_out,
                 Y => Delay1No317_out);

Delay1No318_out_to_Subtract4_0_impl_parent_implementedSystem_port_0_cast <= Delay1No318_out;
Delay1No319_out_to_Subtract4_0_impl_parent_implementedSystem_port_1_cast <= Delay1No319_out;
   Subtract4_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract4_0_impl_out,
                 X => Delay1No318_out_to_Subtract4_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No319_out_to_Subtract4_0_impl_parent_implementedSystem_port_1_cast);

Delay4No210_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_1_cast <= Delay4No210_out;
SharedReg2_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg2_out;
SharedReg646_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg646_out;
SharedReg530_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg530_out;
SharedReg645_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg645_out;
SharedReg645_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg645_out;
SharedReg1006_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1006_out;
SharedReg645_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg645_out;
SharedReg884_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg884_out;
SharedReg127_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg127_out;
SharedReg96_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg96_out;
SharedReg603_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg603_out;
   MUX_Subtract4_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay4No210_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg2_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg96_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg603_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg646_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg530_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg645_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg645_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1006_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg645_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg884_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg127_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract4_0_impl_0_out);

   Delay1No318_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_0_impl_0_out,
                 Y => Delay1No318_out);

SharedReg504_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg504_out;
SharedReg18_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg18_out;
SharedReg822_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg822_out;
SharedReg625_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg625_out;
SharedReg821_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg821_out;
SharedReg821_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg821_out;
SharedReg569_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg569_out;
SharedReg821_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg821_out;
SharedReg961_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg961_out;
SharedReg250_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg250_out;
SharedReg297_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg297_out;
SharedReg645_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg645_out;
   MUX_Subtract4_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg504_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg18_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg297_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg645_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg822_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg625_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg821_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg821_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg569_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg821_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg961_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg250_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract4_0_impl_1_out);

   Delay1No319_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_0_impl_1_out,
                 Y => Delay1No319_out);

Delay1No320_out_to_Subtract4_1_impl_parent_implementedSystem_port_0_cast <= Delay1No320_out;
Delay1No321_out_to_Subtract4_1_impl_parent_implementedSystem_port_1_cast <= Delay1No321_out;
   Subtract4_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract4_1_impl_out,
                 X => Delay1No320_out_to_Subtract4_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No321_out_to_Subtract4_1_impl_parent_implementedSystem_port_1_cast);

SharedReg673_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg673_out;
SharedReg606_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg606_out;
Delay4No211_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_3_cast <= Delay4No211_out;
SharedReg2_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg2_out;
SharedReg649_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg649_out;
SharedReg649_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg649_out;
SharedReg887_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg887_out;
SharedReg887_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg887_out;
SharedReg256_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg256_out;
SharedReg570_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg570_out;
SharedReg779_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg779_out;
SharedReg570_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg570_out;
   MUX_Subtract4_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg673_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg606_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg779_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg570_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => Delay4No211_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg2_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg649_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg649_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg887_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg887_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg256_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg570_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract4_1_impl_0_out);

   Delay1No320_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_1_impl_0_out,
                 Y => Delay1No320_out);

SharedReg672_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg672_out;
SharedReg648_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg648_out;
SharedReg508_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg508_out;
SharedReg18_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg18_out;
SharedReg826_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg826_out;
SharedReg826_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg826_out;
SharedReg963_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg963_out;
SharedReg963_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg963_out;
SharedReg341_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg341_out;
SharedReg854_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg854_out;
SharedReg1007_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1007_out;
SharedReg855_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg855_out;
   MUX_Subtract4_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg672_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg648_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1007_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg855_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg508_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg18_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg826_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg826_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg963_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg963_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg341_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg854_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract4_1_impl_1_out);

   Delay1No321_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_1_impl_1_out,
                 Y => Delay1No321_out);

Delay1No322_out_to_Subtract4_2_impl_parent_implementedSystem_port_0_cast <= Delay1No322_out;
Delay1No323_out_to_Subtract4_2_impl_parent_implementedSystem_port_1_cast <= Delay1No323_out;
   Subtract4_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract4_2_impl_out,
                 X => Delay1No322_out_to_Subtract4_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No323_out_to_Subtract4_2_impl_parent_implementedSystem_port_1_cast);

SharedReg346_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg346_out;
SharedReg445_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg445_out;
SharedReg577_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg577_out;
SharedReg609_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg609_out;
Delay4No212_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_5_cast <= Delay4No212_out;
SharedReg3_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg3_out;
SharedReg946_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg946_out;
SharedReg892_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg892_out;
SharedReg536_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg536_out;
SharedReg1012_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1012_out;
SharedReg1049_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1049_out;
SharedReg879_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg879_out;
   MUX_Subtract4_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg346_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg445_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1049_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg879_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg577_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg609_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay4No212_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg3_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg946_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg892_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg536_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1012_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract4_2_impl_0_out);

   Delay1No322_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_2_impl_0_out,
                 Y => Delay1No322_out);

SharedReg342_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg342_out;
SharedReg679_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg679_out;
SharedReg576_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg576_out;
SharedReg651_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg651_out;
SharedReg512_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg512_out;
SharedReg19_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg19_out;
SharedReg947_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg947_out;
SharedReg967_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg967_out;
SharedReg631_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg631_out;
SharedReg576_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg576_out;
SharedReg449_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg449_out;
SharedReg746_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg746_out;
   MUX_Subtract4_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg342_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg679_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg449_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg746_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg576_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg651_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg512_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg19_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg947_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg967_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg631_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg576_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract4_2_impl_1_out);

   Delay1No323_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_2_impl_1_out,
                 Y => Delay1No323_out);

Delay1No324_out_to_Subtract4_3_impl_parent_implementedSystem_port_0_cast <= Delay1No324_out;
Delay1No325_out_to_Subtract4_3_impl_parent_implementedSystem_port_1_cast <= Delay1No325_out;
   Subtract4_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract4_3_impl_out,
                 X => Delay1No324_out_to_Subtract4_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No325_out_to_Subtract4_3_impl_parent_implementedSystem_port_1_cast);

SharedReg793_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg793_out;
SharedReg455_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg455_out;
SharedReg451_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg451_out;
SharedReg45_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg45_out;
SharedReg612_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg612_out;
Delay4No213_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_6_cast <= Delay4No213_out;
SharedReg2_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg2_out;
SharedReg949_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg949_out;
SharedReg655_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg655_out;
SharedReg539_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg539_out;
SharedReg1017_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1017_out;
SharedReg1055_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1055_out;
   MUX_Subtract4_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg793_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg455_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1017_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1055_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg451_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg45_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg612_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay4No213_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg2_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg949_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg655_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg539_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract4_3_impl_0_out);

   Delay1No324_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_3_impl_0_out,
                 Y => Delay1No324_out);

SharedReg753_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg753_out;
SharedReg1017_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1017_out;
SharedReg862_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg862_out;
SharedReg244_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg244_out;
SharedReg654_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg654_out;
SharedReg516_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg516_out;
SharedReg18_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg18_out;
SharedReg950_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg950_out;
SharedReg834_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg834_out;
SharedReg634_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg634_out;
SharedReg580_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg580_out;
SharedReg457_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg457_out;
   MUX_Subtract4_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg753_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1017_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg580_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg457_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg862_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg244_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg654_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg516_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg18_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg950_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg834_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg634_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract4_3_impl_1_out);

   Delay1No325_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_3_impl_1_out,
                 Y => Delay1No325_out);

Delay1No326_out_to_Subtract4_4_impl_parent_implementedSystem_port_0_cast <= Delay1No326_out;
Delay1No327_out_to_Subtract4_4_impl_parent_implementedSystem_port_1_cast <= Delay1No327_out;
   Subtract4_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract4_4_impl_out,
                 X => Delay1No326_out_to_Subtract4_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No327_out_to_Subtract4_4_impl_parent_implementedSystem_port_1_cast);

SharedReg53_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg53_out;
SharedReg797_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg797_out;
SharedReg767_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg767_out;
SharedReg708_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg708_out;
SharedReg705_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg705_out;
SharedReg459_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg459_out;
SharedReg615_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg615_out;
SharedReg902_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg902_out;
SharedReg3_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg3_out;
SharedReg7_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg7_out;
SharedReg617_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg617_out;
SharedReg658_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg658_out;
   MUX_Subtract4_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg53_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg797_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg617_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg658_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg767_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg708_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg705_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg459_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg615_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg902_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg3_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg7_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract4_4_impl_0_out);

   Delay1No326_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_4_impl_0_out,
                 Y => Delay1No326_out);

SharedReg308_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg308_out;
SharedReg463_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg463_out;
SharedReg758_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg758_out;
SharedReg865_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg865_out;
SharedReg585_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg585_out;
SharedReg458_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg458_out;
SharedReg657_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg657_out;
Delay4No270_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_8_cast <= Delay4No270_out;
SharedReg19_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg19_out;
SharedReg23_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg23_out;
SharedReg902_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg902_out;
SharedReg838_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg838_out;
   MUX_Subtract4_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg308_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg463_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg902_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg838_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg758_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg865_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg585_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg458_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg657_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay4No270_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg19_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg23_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract4_4_impl_1_out);

   Delay1No327_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_4_impl_1_out,
                 Y => Delay1No327_out);

Delay1No328_out_to_Subtract4_5_impl_parent_implementedSystem_port_0_cast <= Delay1No328_out;
Delay1No329_out_to_Subtract4_5_impl_parent_implementedSystem_port_1_cast <= Delay1No329_out;
   Subtract4_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract4_5_impl_out,
                 X => Delay1No328_out_to_Subtract4_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No329_out_to_Subtract4_5_impl_parent_implementedSystem_port_1_cast);

SharedReg620_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg620_out;
SharedReg545_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg545_out;
SharedReg997_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg997_out;
SharedReg292_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg292_out;
SharedReg712_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg712_out;
SharedReg715_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg715_out;
SharedReg150_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg150_out;
SharedReg590_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg590_out;
SharedReg618_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg618_out;
SharedReg906_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg906_out;
SharedReg4_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg7_out;
   MUX_Subtract4_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg620_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg545_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg4_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg7_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg997_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg292_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg712_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg715_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg150_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg590_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg618_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg906_out_to_MUX_Subtract4_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract4_5_impl_0_out);

   Delay1No328_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_5_impl_0_out,
                 Y => Delay1No328_out);

SharedReg906_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg906_out;
SharedReg640_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg640_out;
SharedReg464_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg464_out;
SharedReg319_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg319_out;
SharedReg589_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg589_out;
SharedReg868_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg868_out;
SharedReg183_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg183_out;
SharedReg589_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg589_out;
SharedReg660_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg660_out;
Delay4No271_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_10_cast <= Delay4No271_out;
SharedReg20_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg20_out;
SharedReg23_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg23_out;
   MUX_Subtract4_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg906_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg640_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg20_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg23_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg464_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg319_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg589_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg868_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg183_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg589_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg660_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay4No271_out_to_MUX_Subtract4_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract4_5_impl_1_out);

   Delay1No329_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_5_impl_1_out,
                 Y => Delay1No329_out);

Delay1No330_out_to_Subtract4_6_impl_parent_implementedSystem_port_0_cast <= Delay1No330_out;
Delay1No331_out_to_Subtract4_6_impl_parent_implementedSystem_port_1_cast <= Delay1No331_out;
   Subtract4_6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract4_6_impl_out,
                 X => Delay1No330_out_to_Subtract4_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No331_out_to_Subtract4_6_impl_parent_implementedSystem_port_1_cast);

SharedReg958_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg958_out;
SharedReg548_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg548_out;
SharedReg907_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg907_out;
SharedReg663_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg663_out;
SharedReg1035_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1035_out;
SharedReg663_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg663_out;
SharedReg907_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg907_out;
SharedReg123_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg123_out;
SharedReg771_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg771_out;
SharedReg621_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg621_out;
Delay4No216_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_11_cast <= Delay4No216_out;
SharedReg2_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg2_out;
   MUX_Subtract4_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg958_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg548_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay4No216_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg2_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg907_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg663_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1035_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg663_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg907_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg123_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg771_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg621_out_to_MUX_Subtract4_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract4_6_impl_0_out);

   Delay1No330_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_6_impl_0_out,
                 Y => Delay1No330_out);

SharedReg959_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg959_out;
SharedReg643_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg643_out;
SharedReg978_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg978_out;
SharedReg845_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg845_out;
SharedReg602_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg602_out;
SharedReg845_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg845_out;
SharedReg978_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg978_out;
SharedReg219_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg219_out;
SharedReg595_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg595_out;
SharedReg663_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg663_out;
SharedReg528_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg528_out;
SharedReg18_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg18_out;
   MUX_Subtract4_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg959_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg643_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg528_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg18_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg978_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg845_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg602_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg845_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg978_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg219_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg595_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg663_out_to_MUX_Subtract4_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract4_6_impl_1_out);

   Delay1No331_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_6_impl_1_out,
                 Y => Delay1No331_out);

Delay1No332_out_to_Subtract5_4_impl_parent_implementedSystem_port_0_cast <= Delay1No332_out;
Delay1No333_out_to_Subtract5_4_impl_parent_implementedSystem_port_1_cast <= Delay1No333_out;
   Subtract5_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract5_4_impl_out,
                 X => Delay1No332_out_to_Subtract5_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No333_out_to_Subtract5_4_impl_parent_implementedSystem_port_1_cast);

SharedReg657_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg657_out;
SharedReg541_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg541_out;
SharedReg541_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg541_out;
SharedReg492_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg492_out;
SharedReg616_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg616_out;
SharedReg636_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg636_out;
SharedReg15_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg15_out;
SharedReg424_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg424_out;
SharedReg_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg_out;
SharedReg736_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg736_out;
SharedReg542_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg542_out;
SharedReg657_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg657_out;
   MUX_Subtract5_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg657_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg541_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg542_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg657_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg541_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg492_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg616_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg636_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg15_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg424_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg736_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract5_4_impl_0_out);

   Delay1No332_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract5_4_impl_0_out,
                 Y => Delay1No332_out);

SharedReg837_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg837_out;
SharedReg636_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg636_out;
SharedReg636_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg636_out;
SharedReg558_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg558_out;
SharedReg425_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg425_out;
SharedReg812_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg812_out;
SharedReg31_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg31_out;
SharedReg407_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg407_out;
SharedReg16_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg16_out;
SharedReg559_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg559_out;
SharedReg637_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg637_out;
SharedReg837_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg837_out;
   MUX_Subtract5_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg837_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg636_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg637_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg837_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg636_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg558_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg425_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg812_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg31_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg407_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg16_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg559_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract5_4_impl_1_out);

   Delay1No333_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract5_4_impl_1_out,
                 Y => Delay1No333_out);

Delay1No334_out_to_Subtract5_5_impl_parent_implementedSystem_port_0_cast <= Delay1No334_out;
Delay1No335_out_to_Subtract5_5_impl_parent_implementedSystem_port_1_cast <= Delay1No335_out;
   Subtract5_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract5_5_impl_out,
                 X => Delay1No334_out_to_Subtract5_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No335_out_to_Subtract5_5_impl_parent_implementedSystem_port_1_cast);

SharedReg545_out_to_MUX_Subtract5_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg545_out;
SharedReg544_out_to_MUX_Subtract5_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg544_out;
SharedReg544_out_to_MUX_Subtract5_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg544_out;
SharedReg410_out_to_MUX_Subtract5_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg410_out;
SharedReg410_out_to_MUX_Subtract5_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg410_out;
SharedReg495_out_to_MUX_Subtract5_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg495_out;
SharedReg149_out_to_MUX_Subtract5_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg149_out;
SharedReg639_out_to_MUX_Subtract5_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg639_out;
SharedReg15_out_to_MUX_Subtract5_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg15_out;
SharedReg426_out_to_MUX_Subtract5_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg426_out;
SharedReg1_out_to_MUX_Subtract5_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1_out;
SharedReg740_out_to_MUX_Subtract5_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg740_out;
   MUX_Subtract5_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg545_out_to_MUX_Subtract5_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg544_out_to_MUX_Subtract5_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1_out_to_MUX_Subtract5_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg740_out_to_MUX_Subtract5_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg544_out_to_MUX_Subtract5_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg410_out_to_MUX_Subtract5_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg410_out_to_MUX_Subtract5_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg495_out_to_MUX_Subtract5_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg149_out_to_MUX_Subtract5_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg639_out_to_MUX_Subtract5_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg15_out_to_MUX_Subtract5_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg426_out_to_MUX_Subtract5_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract5_5_impl_0_out);

   Delay1No334_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract5_5_impl_0_out,
                 Y => Delay1No334_out);

SharedReg640_out_to_MUX_Subtract5_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg640_out;
SharedReg639_out_to_MUX_Subtract5_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg639_out;
SharedReg639_out_to_MUX_Subtract5_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg639_out;
SharedReg521_out_to_MUX_Subtract5_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg521_out;
SharedReg521_out_to_MUX_Subtract5_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg521_out;
SharedReg560_out_to_MUX_Subtract5_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg560_out;
SharedReg57_out_to_MUX_Subtract5_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg57_out;
SharedReg815_out_to_MUX_Subtract5_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg815_out;
SharedReg31_out_to_MUX_Subtract5_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg31_out;
SharedReg410_out_to_MUX_Subtract5_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg410_out;
SharedReg17_out_to_MUX_Subtract5_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg17_out;
SharedReg561_out_to_MUX_Subtract5_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg561_out;
   MUX_Subtract5_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg640_out_to_MUX_Subtract5_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg639_out_to_MUX_Subtract5_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg17_out_to_MUX_Subtract5_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg561_out_to_MUX_Subtract5_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg639_out_to_MUX_Subtract5_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg521_out_to_MUX_Subtract5_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg521_out_to_MUX_Subtract5_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg560_out_to_MUX_Subtract5_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg57_out_to_MUX_Subtract5_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg815_out_to_MUX_Subtract5_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg31_out_to_MUX_Subtract5_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg410_out_to_MUX_Subtract5_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract5_5_impl_1_out);

   Delay1No335_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract5_5_impl_1_out,
                 Y => Delay1No335_out);

Delay1No336_out_to_Product26_0_impl_parent_implementedSystem_port_0_cast <= Delay1No336_out;
Delay1No337_out_to_Product26_0_impl_parent_implementedSystem_port_1_cast <= Delay1No337_out;
   Product26_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product26_0_impl_out,
                 X => Delay1No336_out_to_Product26_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No337_out_to_Product26_0_impl_parent_implementedSystem_port_1_cast);

SharedReg1129_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1129_out;
SharedReg1109_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1109_out;
SharedReg1111_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1111_out;
SharedReg1137_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1137_out;
SharedReg1135_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1135_out;
SharedReg1114_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1114_out;
SharedReg1115_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1115_out;
SharedReg1144_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1144_out;
SharedReg1105_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1105_out;
SharedReg1106_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1106_out;
SharedReg1107_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1113_out;
   MUX_Product26_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1129_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1109_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1107_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1113_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1111_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1137_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1135_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1114_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1115_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1144_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1105_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1106_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product26_0_impl_0_out);

   Delay1No336_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product26_0_impl_0_out,
                 Y => Delay1No336_out);

SharedReg1004_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1004_out;
SharedReg1038_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1038_out;
SharedReg127_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg127_out;
SharedReg981_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg981_out;
SharedReg983_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg983_out;
SharedReg1098_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1098_out;
SharedReg202_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg202_out;
SharedReg1071_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1071_out;
SharedReg298_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg298_out;
SharedReg203_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg203_out;
SharedReg1004_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1004_out;
SharedReg1097_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1097_out;
   MUX_Product26_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1004_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1038_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1004_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1097_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg127_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg981_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg983_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1098_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg202_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1071_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg298_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg203_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product26_0_impl_1_out);

   Delay1No337_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product26_0_impl_1_out,
                 Y => Delay1No337_out);

Delay1No338_out_to_Product26_1_impl_parent_implementedSystem_port_0_cast <= Delay1No338_out;
Delay1No339_out_to_Product26_1_impl_parent_implementedSystem_port_1_cast <= Delay1No339_out;
   Product26_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product26_1_impl_out,
                 X => Delay1No338_out_to_Product26_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No339_out_to_Product26_1_impl_parent_implementedSystem_port_1_cast);

SharedReg1107_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1113_out;
SharedReg1129_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1129_out;
SharedReg1109_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1109_out;
SharedReg1111_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1111_out;
SharedReg1137_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1137_out;
SharedReg1135_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1135_out;
SharedReg1114_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1114_out;
SharedReg1115_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1115_out;
SharedReg1144_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1144_out;
SharedReg1105_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1105_out;
SharedReg1106_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1106_out;
   MUX_Product26_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1107_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1113_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1105_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1106_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1129_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1109_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1111_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1137_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1135_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1114_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1115_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1144_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product26_1_impl_0_out);

   Delay1No338_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product26_1_impl_0_out,
                 Y => Delay1No338_out);

SharedReg984_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg984_out;
SharedReg1084_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1084_out;
SharedReg984_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg984_out;
SharedReg1008_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1008_out;
SharedReg100_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg100_out;
SharedReg854_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg854_out;
SharedReg856_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg856_out;
SharedReg1085_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1085_out;
SharedReg234_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg234_out;
SharedReg1082_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1082_out;
SharedReg337_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg337_out;
SharedReg236_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg236_out;
   MUX_Product26_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg984_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1084_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg337_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg236_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg984_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1008_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg100_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg854_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg856_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1085_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg234_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1082_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product26_1_impl_1_out);

   Delay1No339_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product26_1_impl_1_out,
                 Y => Delay1No339_out);

Delay1No340_out_to_Product26_2_impl_parent_implementedSystem_port_0_cast <= Delay1No340_out;
Delay1No341_out_to_Product26_2_impl_parent_implementedSystem_port_1_cast <= Delay1No341_out;
   Product26_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product26_2_impl_out,
                 X => Delay1No340_out_to_Product26_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No341_out_to_Product26_2_impl_parent_implementedSystem_port_1_cast);

SharedReg1105_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1105_out;
SharedReg1106_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1106_out;
SharedReg1107_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1113_out;
SharedReg1129_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1129_out;
SharedReg1109_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1109_out;
SharedReg1111_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1111_out;
SharedReg1137_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1137_out;
SharedReg1135_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1135_out;
SharedReg1114_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1114_out;
SharedReg1115_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1115_out;
SharedReg1144_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1144_out;
   MUX_Product26_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1105_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1106_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1115_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1144_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1107_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1113_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1129_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1109_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1111_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1137_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1135_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1114_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product26_2_impl_0_out);

   Delay1No340_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product26_2_impl_0_out,
                 Y => Delay1No340_out);

SharedReg304_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg304_out;
SharedReg241_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg241_out;
SharedReg858_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg858_out;
SharedReg1050_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1050_out;
SharedReg858_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg858_out;
SharedReg987_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg987_out;
SharedReg134_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg134_out;
SharedReg858_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg858_out;
SharedReg680_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg680_out;
SharedReg1051_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1051_out;
SharedReg239_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg239_out;
SharedReg1048_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1048_out;
   MUX_Product26_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg304_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg241_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg239_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1048_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg858_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1050_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg858_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg987_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg134_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg858_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg680_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1051_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product26_2_impl_1_out);

   Delay1No341_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product26_2_impl_1_out,
                 Y => Delay1No341_out);

Delay1No342_out_to_Product26_3_impl_parent_implementedSystem_port_0_cast <= Delay1No342_out;
Delay1No343_out_to_Product26_3_impl_parent_implementedSystem_port_1_cast <= Delay1No343_out;
   Product26_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product26_3_impl_out,
                 X => Delay1No342_out_to_Product26_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No343_out_to_Product26_3_impl_parent_implementedSystem_port_1_cast);

SharedReg1144_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1144_out;
SharedReg1105_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1105_out;
SharedReg1106_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1106_out;
SharedReg1107_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1113_out;
SharedReg1129_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1129_out;
SharedReg1109_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1109_out;
SharedReg1111_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1111_out;
SharedReg1137_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1137_out;
SharedReg1135_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1135_out;
SharedReg1114_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1114_out;
SharedReg1115_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1115_out;
   MUX_Product26_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1144_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1105_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1114_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1115_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1106_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1107_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1113_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1129_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1109_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1111_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1137_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1135_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product26_3_impl_0_out);

   Delay1No342_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product26_3_impl_0_out,
                 Y => Delay1No342_out);

SharedReg791_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg791_out;
SharedReg352_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg352_out;
SharedReg141_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg141_out;
SharedReg861_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg861_out;
SharedReg793_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg793_out;
SharedReg861_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg861_out;
SharedReg991_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg991_out;
SharedReg110_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg110_out;
SharedReg990_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg990_out;
SharedReg863_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg863_out;
SharedReg1057_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1057_out;
SharedReg244_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg244_out;
   MUX_Product26_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg791_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg352_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1057_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg244_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg141_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg861_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg793_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg861_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg991_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg110_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg990_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg863_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product26_3_impl_1_out);

   Delay1No343_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product26_3_impl_1_out,
                 Y => Delay1No343_out);

Delay1No344_out_to_Product26_4_impl_parent_implementedSystem_port_0_cast <= Delay1No344_out;
Delay1No345_out_to_Product26_4_impl_parent_implementedSystem_port_1_cast <= Delay1No345_out;
   Product26_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product26_4_impl_out,
                 X => Delay1No344_out_to_Product26_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No345_out_to_Product26_4_impl_parent_implementedSystem_port_1_cast);

SharedReg1114_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1114_out;
SharedReg1115_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1115_out;
SharedReg1144_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1144_out;
SharedReg1105_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1105_out;
SharedReg1106_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1106_out;
SharedReg1107_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1113_out;
SharedReg1129_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1129_out;
SharedReg1109_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1109_out;
SharedReg1111_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1111_out;
SharedReg1137_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1137_out;
SharedReg1135_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1135_out;
   MUX_Product26_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1114_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1115_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1137_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1135_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1144_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1105_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1106_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1107_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1113_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1129_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1109_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1111_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product26_4_impl_0_out);

   Delay1No344_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product26_4_impl_0_out,
                 Y => Delay1No344_out);

SharedReg799_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg799_out;
SharedReg206_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg206_out;
SharedReg796_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg796_out;
SharedReg310_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg310_out;
SharedReg147_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg147_out;
SharedReg689_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg689_out;
SharedReg1024_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1024_out;
SharedReg865_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg865_out;
SharedReg994_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg994_out;
SharedReg145_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg145_out;
SharedReg865_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg865_out;
SharedReg867_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg867_out;
   MUX_Product26_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg799_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg206_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg865_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg867_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg796_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg310_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg147_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg689_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1024_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg865_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg994_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg145_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product26_4_impl_1_out);

   Delay1No345_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product26_4_impl_1_out,
                 Y => Delay1No345_out);

Delay1No346_out_to_Product26_5_impl_parent_implementedSystem_port_0_cast <= Delay1No346_out;
Delay1No347_out_to_Product26_5_impl_parent_implementedSystem_port_1_cast <= Delay1No347_out;
   Product26_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product26_5_impl_out,
                 X => Delay1No346_out_to_Product26_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No347_out_to_Product26_5_impl_parent_implementedSystem_port_1_cast);

SharedReg1137_out_to_MUX_Product26_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1137_out;
SharedReg1135_out_to_MUX_Product26_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1135_out;
SharedReg1114_out_to_MUX_Product26_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1114_out;
SharedReg1115_out_to_MUX_Product26_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1115_out;
SharedReg1144_out_to_MUX_Product26_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1144_out;
SharedReg1105_out_to_MUX_Product26_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1105_out;
SharedReg1106_out_to_MUX_Product26_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1106_out;
SharedReg1107_out_to_MUX_Product26_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product26_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1113_out;
SharedReg1129_out_to_MUX_Product26_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1129_out;
SharedReg1109_out_to_MUX_Product26_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1109_out;
SharedReg1111_out_to_MUX_Product26_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1111_out;
   MUX_Product26_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1137_out_to_MUX_Product26_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1135_out_to_MUX_Product26_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1109_out_to_MUX_Product26_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1111_out_to_MUX_Product26_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1114_out_to_MUX_Product26_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1115_out_to_MUX_Product26_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1144_out_to_MUX_Product26_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1105_out_to_MUX_Product26_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1106_out_to_MUX_Product26_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1107_out_to_MUX_Product26_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1113_out_to_MUX_Product26_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1129_out_to_MUX_Product26_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product26_5_impl_0_out);

   Delay1No346_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product26_5_impl_0_out,
                 Y => Delay1No346_out);

SharedReg868_out_to_MUX_Product26_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg868_out;
SharedReg870_out_to_MUX_Product26_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg870_out;
SharedReg774_out_to_MUX_Product26_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg774_out;
SharedReg182_out_to_MUX_Product26_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg182_out;
SharedReg1029_out_to_MUX_Product26_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1029_out;
SharedReg288_out_to_MUX_Product26_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg288_out;
SharedReg184_out_to_MUX_Product26_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg184_out;
SharedReg868_out_to_MUX_Product26_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg868_out;
SharedReg1031_out_to_MUX_Product26_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1031_out;
SharedReg997_out_to_MUX_Product26_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg997_out;
SharedReg1029_out_to_MUX_Product26_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1029_out;
SharedReg212_out_to_MUX_Product26_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg212_out;
   MUX_Product26_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg868_out_to_MUX_Product26_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg870_out_to_MUX_Product26_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1029_out_to_MUX_Product26_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg212_out_to_MUX_Product26_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg774_out_to_MUX_Product26_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg182_out_to_MUX_Product26_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1029_out_to_MUX_Product26_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg288_out_to_MUX_Product26_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg184_out_to_MUX_Product26_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg868_out_to_MUX_Product26_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1031_out_to_MUX_Product26_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg997_out_to_MUX_Product26_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product26_5_impl_1_out);

   Delay1No347_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product26_5_impl_1_out,
                 Y => Delay1No347_out);

Delay1No348_out_to_Product26_6_impl_parent_implementedSystem_port_0_cast <= Delay1No348_out;
Delay1No349_out_to_Product26_6_impl_parent_implementedSystem_port_1_cast <= Delay1No349_out;
   Product26_6_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product26_6_impl_out,
                 X => Delay1No348_out_to_Product26_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No349_out_to_Product26_6_impl_parent_implementedSystem_port_1_cast);

SharedReg1111_out_to_MUX_Product26_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1111_out;
SharedReg1137_out_to_MUX_Product26_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1137_out;
SharedReg1135_out_to_MUX_Product26_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1135_out;
SharedReg1114_out_to_MUX_Product26_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1114_out;
SharedReg1115_out_to_MUX_Product26_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1115_out;
SharedReg1144_out_to_MUX_Product26_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1144_out;
SharedReg1105_out_to_MUX_Product26_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1105_out;
SharedReg1106_out_to_MUX_Product26_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1106_out;
SharedReg1107_out_to_MUX_Product26_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1107_out;
SharedReg1113_out_to_MUX_Product26_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1113_out;
SharedReg1129_out_to_MUX_Product26_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1129_out;
SharedReg1109_out_to_MUX_Product26_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1109_out;
   MUX_Product26_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1111_out_to_MUX_Product26_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1137_out_to_MUX_Product26_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1129_out_to_MUX_Product26_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1109_out_to_MUX_Product26_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1135_out_to_MUX_Product26_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1114_out_to_MUX_Product26_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1115_out_to_MUX_Product26_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1144_out_to_MUX_Product26_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1105_out_to_MUX_Product26_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1106_out_to_MUX_Product26_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1107_out_to_MUX_Product26_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1113_out_to_MUX_Product26_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product26_6_impl_0_out);

   Delay1No348_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product26_6_impl_0_out,
                 Y => Delay1No348_out);

SharedReg153_out_to_MUX_Product26_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg153_out;
SharedReg1033_out_to_MUX_Product26_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1033_out;
SharedReg1036_out_to_MUX_Product26_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1036_out;
SharedReg1092_out_to_MUX_Product26_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1092_out;
SharedReg187_out_to_MUX_Product26_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg187_out;
SharedReg1076_out_to_MUX_Product26_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1076_out;
SharedReg322_out_to_MUX_Product26_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg322_out;
SharedReg155_out_to_MUX_Product26_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg155_out;
SharedReg1033_out_to_MUX_Product26_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1033_out;
SharedReg1091_out_to_MUX_Product26_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1091_out;
SharedReg1033_out_to_MUX_Product26_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1033_out;
SharedReg1067_out_to_MUX_Product26_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1067_out;
   MUX_Product26_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg153_out_to_MUX_Product26_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1033_out_to_MUX_Product26_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1033_out_to_MUX_Product26_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1067_out_to_MUX_Product26_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1036_out_to_MUX_Product26_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1092_out_to_MUX_Product26_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg187_out_to_MUX_Product26_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1076_out_to_MUX_Product26_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg322_out_to_MUX_Product26_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg155_out_to_MUX_Product26_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1033_out_to_MUX_Product26_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1091_out_to_MUX_Product26_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product26_6_impl_1_out);

   Delay1No349_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product26_6_impl_1_out,
                 Y => Delay1No349_out);

Delay1No350_out_to_Subtract7_2_impl_parent_implementedSystem_port_0_cast <= Delay1No350_out;
Delay1No351_out_to_Subtract7_2_impl_parent_implementedSystem_port_1_cast <= Delay1No351_out;
   Subtract7_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract7_2_impl_out,
                 X => Delay1No350_out_to_Subtract7_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No351_out_to_Subtract7_2_impl_parent_implementedSystem_port_1_cast);

SharedReg891_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg891_out;
SharedReg610_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg610_out;
SharedReg630_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg630_out;
SharedReg15_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg15_out;
SharedReg14_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg14_out;
SharedReg_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg_out;
SharedReg653_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg653_out;
SharedReg402_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg402_out;
SharedReg535_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg535_out;
SharedReg535_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg535_out;
SharedReg535_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg535_out;
SharedReg535_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg535_out;
   MUX_Subtract7_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg891_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg610_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg535_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg535_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg630_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg15_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg14_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg653_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg402_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg535_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg535_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract7_2_impl_0_out);

   Delay1No350_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract7_2_impl_0_out,
                 Y => Delay1No350_out);

SharedReg966_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg966_out;
SharedReg421_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg421_out;
SharedReg806_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg806_out;
SharedReg31_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg31_out;
SharedReg30_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg30_out;
SharedReg16_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg16_out;
SharedReg421_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg421_out;
SharedReg510_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg510_out;
SharedReg630_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg630_out;
SharedReg630_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg630_out;
SharedReg630_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg630_out;
SharedReg630_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg630_out;
   MUX_Subtract7_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg966_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg421_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg630_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg630_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg806_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg31_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg30_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg16_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg421_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg510_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg630_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg630_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract7_2_impl_1_out);

   Delay1No351_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract7_2_impl_1_out,
                 Y => Delay1No351_out);

Delay1No352_out_to_Subtract7_3_impl_parent_implementedSystem_port_0_cast <= Delay1No352_out;
Delay1No353_out_to_Subtract7_3_impl_parent_implementedSystem_port_1_cast <= Delay1No353_out;
   Subtract7_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract7_3_impl_out,
                 X => Delay1No352_out_to_Subtract7_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No353_out_to_Subtract7_3_impl_parent_implementedSystem_port_1_cast);

SharedReg538_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg538_out;
SharedReg489_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg489_out;
SharedReg613_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg613_out;
SharedReg243_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg243_out;
SharedReg860_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg860_out;
SharedReg15_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg15_out;
SharedReg14_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg14_out;
SharedReg656_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg656_out;
SharedReg491_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg491_out;
SharedReg538_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg538_out;
SharedReg538_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg538_out;
SharedReg538_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg538_out;
   MUX_Subtract7_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg538_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg489_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg538_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg538_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg613_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg243_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg860_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg15_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg14_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg656_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg491_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg538_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract7_3_impl_0_out);

   Delay1No352_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract7_3_impl_0_out,
                 Y => Delay1No352_out);

SharedReg633_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg633_out;
SharedReg556_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg556_out;
SharedReg423_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg423_out;
SharedReg174_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg174_out;
SharedReg450_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg450_out;
SharedReg31_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg31_out;
SharedReg30_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg30_out;
SharedReg423_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg423_out;
Delay6No10_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_9_cast <= Delay6No10_out;
SharedReg633_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg633_out;
SharedReg633_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg633_out;
SharedReg633_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg633_out;
   MUX_Subtract7_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg633_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg556_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg633_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg633_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg423_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg174_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg450_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg31_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg30_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg423_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay6No10_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg633_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract7_3_impl_1_out);

   Delay1No353_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract7_3_impl_1_out,
                 Y => Delay1No353_out);

Delay1No354_out_to_Subtract7_4_impl_parent_implementedSystem_port_0_cast <= Delay1No354_out;
Delay1No355_out_to_Subtract7_4_impl_parent_implementedSystem_port_1_cast <= Delay1No355_out;
   Subtract7_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract7_4_impl_out,
                 X => Delay1No354_out_to_Subtract7_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No355_out_to_Subtract7_4_impl_parent_implementedSystem_port_1_cast);

SharedReg541_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg541_out;
SharedReg407_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg407_out;
SharedReg407_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg407_out;
SharedReg192_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg192_out;
SharedReg144_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg144_out;
SharedReg864_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg864_out;
SharedReg13_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg13_out;
SharedReg14_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg14_out;
SharedReg268_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg268_out;
SharedReg659_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg659_out;
SharedReg408_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg408_out;
SharedReg541_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg541_out;
   MUX_Subtract7_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg541_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg407_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg408_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg541_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg407_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg192_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg144_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg864_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg13_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg14_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg268_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg659_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract7_4_impl_0_out);

   Delay1No354_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract7_4_impl_0_out,
                 Y => Delay1No354_out);

SharedReg636_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg636_out;
SharedReg517_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg517_out;
SharedReg517_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg517_out;
SharedReg353_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg353_out;
SharedReg181_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg181_out;
SharedReg583_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg583_out;
SharedReg29_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg30_out;
SharedReg352_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg352_out;
SharedReg425_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg425_out;
SharedReg518_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg518_out;
SharedReg636_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg636_out;
   MUX_Subtract7_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg636_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg517_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg518_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg636_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg517_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg353_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg181_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg583_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg29_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg30_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg352_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg425_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract7_4_impl_1_out);

   Delay1No355_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract7_4_impl_1_out,
                 Y => Delay1No355_out);

Delay1No356_out_to_Subtract7_5_impl_parent_implementedSystem_port_0_cast <= Delay1No356_out;
Delay1No357_out_to_Subtract7_5_impl_parent_implementedSystem_port_1_cast <= Delay1No357_out;
   Subtract7_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract7_5_impl_out,
                 X => Delay1No356_out_to_Subtract7_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No357_out_to_Subtract7_5_impl_parent_implementedSystem_port_1_cast);

SharedReg411_out_to_MUX_Subtract7_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg411_out;
SharedReg410_out_to_MUX_Subtract7_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg410_out;
SharedReg410_out_to_MUX_Subtract7_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg410_out;
SharedReg461_out_to_MUX_Subtract7_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg461_out;
SharedReg272_out_to_MUX_Subtract7_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg272_out;
SharedReg279_out_to_MUX_Subtract7_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg279_out;
SharedReg952_out_to_MUX_Subtract7_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg952_out;
SharedReg693_out_to_MUX_Subtract7_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg693_out;
SharedReg13_out_to_MUX_Subtract7_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg13_out;
SharedReg14_out_to_MUX_Subtract7_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg14_out;
SharedReg_out_to_MUX_Subtract7_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg_out;
SharedReg662_out_to_MUX_Subtract7_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg662_out;
   MUX_Subtract7_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg411_out_to_MUX_Subtract7_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg410_out_to_MUX_Subtract7_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg_out_to_MUX_Subtract7_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg662_out_to_MUX_Subtract7_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg410_out_to_MUX_Subtract7_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg461_out_to_MUX_Subtract7_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg272_out_to_MUX_Subtract7_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg279_out_to_MUX_Subtract7_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg952_out_to_MUX_Subtract7_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg693_out_to_MUX_Subtract7_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg13_out_to_MUX_Subtract7_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg14_out_to_MUX_Subtract7_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract7_5_impl_0_out);

   Delay1No356_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract7_5_impl_0_out,
                 Y => Delay1No356_out);

SharedReg522_out_to_MUX_Subtract7_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg522_out;
SharedReg521_out_to_MUX_Subtract7_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg521_out;
SharedReg521_out_to_MUX_Subtract7_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg521_out;
SharedReg689_out_to_MUX_Subtract7_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg689_out;
SharedReg276_out_to_MUX_Subtract7_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg276_out;
SharedReg284_out_to_MUX_Subtract7_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg284_out;
SharedReg972_out_to_MUX_Subtract7_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg972_out;
SharedReg588_out_to_MUX_Subtract7_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg588_out;
SharedReg29_out_to_MUX_Subtract7_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Subtract7_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg30_out;
SharedReg16_out_to_MUX_Subtract7_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg16_out;
SharedReg427_out_to_MUX_Subtract7_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg427_out;
   MUX_Subtract7_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg522_out_to_MUX_Subtract7_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg521_out_to_MUX_Subtract7_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg16_out_to_MUX_Subtract7_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg427_out_to_MUX_Subtract7_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg521_out_to_MUX_Subtract7_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg689_out_to_MUX_Subtract7_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg276_out_to_MUX_Subtract7_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg284_out_to_MUX_Subtract7_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg972_out_to_MUX_Subtract7_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg588_out_to_MUX_Subtract7_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg29_out_to_MUX_Subtract7_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg30_out_to_MUX_Subtract7_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract7_5_impl_1_out);

   Delay1No357_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract7_5_impl_1_out,
                 Y => Delay1No357_out);

Delay1No358_out_to_Subtract7_6_impl_parent_implementedSystem_port_0_cast <= Delay1No358_out;
Delay1No359_out_to_Subtract7_6_impl_parent_implementedSystem_port_1_cast <= Delay1No359_out;
   Subtract7_6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract7_6_impl_out,
                 X => Delay1No358_out_to_Subtract7_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No359_out_to_Subtract7_6_impl_parent_implementedSystem_port_1_cast);

SharedReg665_out_to_MUX_Subtract7_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg665_out;
SharedReg470_out_to_MUX_Subtract7_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg470_out;
SharedReg413_out_to_MUX_Subtract7_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg413_out;
SharedReg294_out_to_MUX_Subtract7_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg294_out;
SharedReg152_out_to_MUX_Subtract7_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg152_out;
SharedReg468_out_to_MUX_Subtract7_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg468_out;
SharedReg868_out_to_MUX_Subtract7_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg868_out;
SharedReg225_out_to_MUX_Subtract7_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg225_out;
SharedReg955_out_to_MUX_Subtract7_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg955_out;
SharedReg698_out_to_MUX_Subtract7_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg698_out;
SharedReg15_out_to_MUX_Subtract7_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg15_out;
SharedReg14_out_to_MUX_Subtract7_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg14_out;
   MUX_Subtract7_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg665_out_to_MUX_Subtract7_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg470_out_to_MUX_Subtract7_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg15_out_to_MUX_Subtract7_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg14_out_to_MUX_Subtract7_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg413_out_to_MUX_Subtract7_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg294_out_to_MUX_Subtract7_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg152_out_to_MUX_Subtract7_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg468_out_to_MUX_Subtract7_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg868_out_to_MUX_Subtract7_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg225_out_to_MUX_Subtract7_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg955_out_to_MUX_Subtract7_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg698_out_to_MUX_Subtract7_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract7_6_impl_0_out);

   Delay1No358_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract7_6_impl_0_out,
                 Y => Delay1No358_out);

SharedReg429_out_to_MUX_Subtract7_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg429_out;
SharedReg467_out_to_MUX_Subtract7_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg467_out;
SharedReg525_out_to_MUX_Subtract7_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg525_out;
SharedReg288_out_to_MUX_Subtract7_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg288_out;
SharedReg224_out_to_MUX_Subtract7_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg224_out;
SharedReg694_out_to_MUX_Subtract7_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg694_out;
SharedReg471_out_to_MUX_Subtract7_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg471_out;
SharedReg231_out_to_MUX_Subtract7_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg231_out;
SharedReg975_out_to_MUX_Subtract7_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg975_out;
SharedReg594_out_to_MUX_Subtract7_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg594_out;
SharedReg31_out_to_MUX_Subtract7_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg31_out;
SharedReg30_out_to_MUX_Subtract7_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg30_out;
   MUX_Subtract7_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg429_out_to_MUX_Subtract7_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg467_out_to_MUX_Subtract7_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg31_out_to_MUX_Subtract7_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg30_out_to_MUX_Subtract7_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg525_out_to_MUX_Subtract7_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg288_out_to_MUX_Subtract7_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg224_out_to_MUX_Subtract7_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg694_out_to_MUX_Subtract7_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg471_out_to_MUX_Subtract7_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg231_out_to_MUX_Subtract7_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg975_out_to_MUX_Subtract7_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg594_out_to_MUX_Subtract7_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract7_6_impl_1_out);

   Delay1No359_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract7_6_impl_1_out,
                 Y => Delay1No359_out);

Delay1No360_out_to_Subtract8_1_impl_parent_implementedSystem_port_0_cast <= Delay1No360_out;
Delay1No361_out_to_Subtract8_1_impl_parent_implementedSystem_port_1_cast <= Delay1No361_out;
   Subtract8_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract8_1_impl_out,
                 X => Delay1No360_out_to_Subtract8_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No361_out_to_Subtract8_1_impl_parent_implementedSystem_port_1_cast);

SharedReg627_out_to_MUX_Subtract8_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg627_out;
SharedReg15_out_to_MUX_Subtract8_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg15_out;
SharedReg14_out_to_MUX_Subtract8_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg14_out;
SharedReg299_out_to_MUX_Subtract8_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg299_out;
SharedReg853_out_to_MUX_Subtract8_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg853_out;
SharedReg485_out_to_MUX_Subtract8_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg485_out;
SharedReg398_out_to_MUX_Subtract8_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg398_out;
SharedReg398_out_to_MUX_Subtract8_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg398_out;
SharedReg398_out_to_MUX_Subtract8_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg398_out;
SharedReg398_out_to_MUX_Subtract8_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg398_out;
SharedReg483_out_to_MUX_Subtract8_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg483_out;
SharedReg607_out_to_MUX_Subtract8_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg607_out;
   MUX_Subtract8_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg627_out_to_MUX_Subtract8_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg15_out_to_MUX_Subtract8_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg483_out_to_MUX_Subtract8_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg607_out_to_MUX_Subtract8_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg14_out_to_MUX_Subtract8_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg299_out_to_MUX_Subtract8_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg853_out_to_MUX_Subtract8_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg485_out_to_MUX_Subtract8_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg398_out_to_MUX_Subtract8_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg398_out_to_MUX_Subtract8_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg398_out_to_MUX_Subtract8_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg398_out_to_MUX_Subtract8_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract8_1_impl_0_out);

   Delay1No360_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract8_1_impl_0_out,
                 Y => Delay1No360_out);

SharedReg803_out_to_MUX_Subtract8_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg803_out;
SharedReg31_out_to_MUX_Subtract8_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg31_out;
SharedReg30_out_to_MUX_Subtract8_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg30_out;
SharedReg328_out_to_MUX_Subtract8_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg328_out;
SharedReg566_out_to_MUX_Subtract8_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg566_out;
Delay6No8_out_to_MUX_Subtract8_1_impl_1_parent_implementedSystem_port_6_cast <= Delay6No8_out;
SharedReg505_out_to_MUX_Subtract8_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg505_out;
SharedReg505_out_to_MUX_Subtract8_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg505_out;
SharedReg505_out_to_MUX_Subtract8_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg505_out;
SharedReg505_out_to_MUX_Subtract8_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg505_out;
SharedReg552_out_to_MUX_Subtract8_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg552_out;
SharedReg419_out_to_MUX_Subtract8_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg419_out;
   MUX_Subtract8_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg803_out_to_MUX_Subtract8_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg31_out_to_MUX_Subtract8_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg552_out_to_MUX_Subtract8_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg419_out_to_MUX_Subtract8_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg30_out_to_MUX_Subtract8_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg328_out_to_MUX_Subtract8_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg566_out_to_MUX_Subtract8_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay6No8_out_to_MUX_Subtract8_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg505_out_to_MUX_Subtract8_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg505_out_to_MUX_Subtract8_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg505_out_to_MUX_Subtract8_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg505_out_to_MUX_Subtract8_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract8_1_impl_1_out);

   Delay1No361_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract8_1_impl_1_out,
                 Y => Delay1No361_out);

Delay1No362_out_to_Subtract8_2_impl_parent_implementedSystem_port_0_cast <= Delay1No362_out;
Delay1No363_out_to_Subtract8_2_impl_parent_implementedSystem_port_1_cast <= Delay1No363_out;
   Subtract8_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract8_2_impl_out,
                 X => Delay1No362_out_to_Subtract8_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No363_out_to_Subtract8_2_impl_parent_implementedSystem_port_1_cast);

SharedReg486_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg486_out;
SharedReg238_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg238_out;
SharedReg857_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg857_out;
SharedReg13_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg13_out;
SharedReg12_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg12_out;
SharedReg257_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg257_out;
SharedReg677_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg677_out;
SharedReg488_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg488_out;
SharedReg401_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg401_out;
SharedReg401_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg401_out;
SharedReg401_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg401_out;
SharedReg401_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg401_out;
   MUX_Subtract8_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg486_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg238_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg401_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg401_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg857_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg13_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg12_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg257_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg677_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg488_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg401_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg401_out_to_MUX_Subtract8_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract8_2_impl_0_out);

   Delay1No362_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract8_2_impl_0_out,
                 Y => Delay1No362_out);

SharedReg554_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg554_out;
SharedReg376_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg376_out;
SharedReg575_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg575_out;
SharedReg29_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg29_out;
SharedReg28_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg28_out;
SharedReg337_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg337_out;
SharedReg440_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg440_out;
Delay6No9_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_8_cast <= Delay6No9_out;
SharedReg509_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg509_out;
SharedReg509_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg509_out;
SharedReg509_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg509_out;
SharedReg509_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg509_out;
   MUX_Subtract8_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg554_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg376_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg509_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg509_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg575_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg29_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg28_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg337_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg440_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay6No9_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg509_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg509_out_to_MUX_Subtract8_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract8_2_impl_1_out);

   Delay1No363_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract8_2_impl_1_out,
                 Y => Delay1No363_out);

Delay1No364_out_to_Subtract8_4_impl_parent_implementedSystem_port_0_cast <= Delay1No364_out;
Delay1No365_out_to_Subtract8_4_impl_parent_implementedSystem_port_1_cast <= Delay1No365_out;
   Subtract8_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract8_4_impl_out,
                 X => Delay1No364_out_to_Subtract8_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No365_out_to_Subtract8_4_impl_parent_implementedSystem_port_1_cast);

SharedReg407_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg407_out;
SharedReg454_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg454_out;
SharedReg266_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg266_out;
SharedReg1018_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1018_out;
SharedReg949_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg949_out;
SharedReg195_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg195_out;
SharedReg10_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg10_out;
SharedReg12_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg12_out;
SharedReg113_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg113_out;
SharedReg688_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg688_out;
SharedReg494_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg494_out;
SharedReg407_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg407_out;
   MUX_Subtract8_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg407_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg454_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg494_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg407_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg266_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1018_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg949_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg195_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg10_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg12_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg113_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg688_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract8_4_impl_0_out);

   Delay1No364_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract8_4_impl_0_out,
                 Y => Delay1No364_out);

SharedReg517_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg517_out;
SharedReg990_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg990_out;
SharedReg247_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg247_out;
SharedReg1021_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1021_out;
SharedReg969_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg969_out;
SharedReg248_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg248_out;
SharedReg26_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg26_out;
SharedReg28_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg28_out;
SharedReg267_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg267_out;
SharedReg453_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg453_out;
Delay6No11_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_11_cast <= Delay6No11_out;
SharedReg517_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg517_out;
   MUX_Subtract8_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg517_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg990_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay6No11_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg517_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg247_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1021_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg969_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg248_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg26_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg28_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg267_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg453_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract8_4_impl_1_out);

   Delay1No365_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract8_4_impl_1_out,
                 Y => Delay1No365_out);

Delay1No366_out_to_Subtract8_5_impl_parent_implementedSystem_port_0_cast <= Delay1No366_out;
Delay1No367_out_to_Subtract8_5_impl_parent_implementedSystem_port_1_cast <= Delay1No367_out;
   Subtract8_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract8_5_impl_out,
                 X => Delay1No366_out_to_Subtract8_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No367_out_to_Subtract8_5_impl_parent_implementedSystem_port_1_cast);

SharedReg497_out_to_MUX_Subtract8_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg497_out;
SharedReg275_out_to_MUX_Subtract8_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg275_out;
SharedReg116_out_to_MUX_Subtract8_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg116_out;
SharedReg148_out_to_MUX_Subtract8_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg148_out;
SharedReg689_out_to_MUX_Subtract8_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg689_out;
SharedReg994_out_to_MUX_Subtract8_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg994_out;
SharedReg659_out_to_MUX_Subtract8_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg659_out;
SharedReg283_out_to_MUX_Subtract8_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg283_out;
SharedReg10_out_to_MUX_Subtract8_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg10_out;
SharedReg12_out_to_MUX_Subtract8_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg12_out;
SharedReg210_out_to_MUX_Subtract8_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg210_out;
SharedReg462_out_to_MUX_Subtract8_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg462_out;
   MUX_Subtract8_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg497_out_to_MUX_Subtract8_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg275_out_to_MUX_Subtract8_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg210_out_to_MUX_Subtract8_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg462_out_to_MUX_Subtract8_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg116_out_to_MUX_Subtract8_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg148_out_to_MUX_Subtract8_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg689_out_to_MUX_Subtract8_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg994_out_to_MUX_Subtract8_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg659_out_to_MUX_Subtract8_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg283_out_to_MUX_Subtract8_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg10_out_to_MUX_Subtract8_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg12_out_to_MUX_Subtract8_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract8_5_impl_0_out);

   Delay1No366_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract8_5_impl_0_out,
                 Y => Delay1No366_out);

Delay6No12_out_to_MUX_Subtract8_5_impl_1_parent_implementedSystem_port_1_cast <= Delay6No12_out;
SharedReg274_out_to_MUX_Subtract8_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg274_out;
SharedReg52_out_to_MUX_Subtract8_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg52_out;
SharedReg114_out_to_MUX_Subtract8_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg114_out;
SharedReg710_out_to_MUX_Subtract8_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg710_out;
SharedReg1027_out_to_MUX_Subtract8_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1027_out;
SharedReg839_out_to_MUX_Subtract8_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg839_out;
SharedReg277_out_to_MUX_Subtract8_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg277_out;
SharedReg26_out_to_MUX_Subtract8_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg26_out;
SharedReg28_out_to_MUX_Subtract8_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg28_out;
SharedReg280_out_to_MUX_Subtract8_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg280_out;
SharedReg460_out_to_MUX_Subtract8_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg460_out;
   MUX_Subtract8_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay6No12_out_to_MUX_Subtract8_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg274_out_to_MUX_Subtract8_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg280_out_to_MUX_Subtract8_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg460_out_to_MUX_Subtract8_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg52_out_to_MUX_Subtract8_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg114_out_to_MUX_Subtract8_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg710_out_to_MUX_Subtract8_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1027_out_to_MUX_Subtract8_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg839_out_to_MUX_Subtract8_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg277_out_to_MUX_Subtract8_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg26_out_to_MUX_Subtract8_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg28_out_to_MUX_Subtract8_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract8_5_impl_1_out);

   Delay1No367_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract8_5_impl_1_out,
                 Y => Delay1No367_out);

Delay1No368_out_to_Product18_0_impl_parent_implementedSystem_port_0_cast <= Delay1No368_out;
Delay1No369_out_to_Product18_0_impl_parent_implementedSystem_port_1_cast <= Delay1No369_out;
   Product18_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product18_0_impl_out,
                 X => Delay1No368_out_to_Product18_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No369_out_to_Product18_0_impl_parent_implementedSystem_port_1_cast);

SharedReg1131_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1131_out;
SharedReg1121_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1121_out;
SharedReg1123_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1123_out;
SharedReg1141_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1141_out;
SharedReg1139_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1139_out;
SharedReg1126_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1126_out;
SharedReg249_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg249_out;
SharedReg1155_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1155_out;
SharedReg1117_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1117_out;
SharedReg1118_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1118_out;
SharedReg1119_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1125_out;
   MUX_Product18_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1131_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1121_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1119_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1125_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1123_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1141_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1139_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1126_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg249_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1155_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1117_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1118_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product18_0_impl_0_out);

   Delay1No368_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product18_0_impl_0_out,
                 Y => Delay1No368_out);

SharedReg981_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg981_out;
SharedReg1094_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1094_out;
SharedReg32_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg32_out;
SharedReg849_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg849_out;
SharedReg851_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg851_out;
SharedReg1099_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1099_out;
SharedReg1115_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1115_out;
SharedReg775_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg775_out;
SharedReg298_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg298_out;
SharedReg329_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg329_out;
SharedReg981_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg981_out;
SharedReg1073_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1073_out;
   MUX_Product18_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg981_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1094_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg981_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1073_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg32_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg849_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg851_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1099_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1115_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg775_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg298_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg329_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product18_0_impl_1_out);

   Delay1No369_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product18_0_impl_1_out,
                 Y => Delay1No369_out);

Delay1No370_out_to_Product18_1_impl_parent_implementedSystem_port_0_cast <= Delay1No370_out;
Delay1No371_out_to_Product18_1_impl_parent_implementedSystem_port_1_cast <= Delay1No371_out;
   Product18_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product18_1_impl_out,
                 X => Delay1No370_out_to_Product18_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No371_out_to_Product18_1_impl_parent_implementedSystem_port_1_cast);

SharedReg1119_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1125_out;
SharedReg1131_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1131_out;
SharedReg1121_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1121_out;
SharedReg1123_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1123_out;
SharedReg1141_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1141_out;
SharedReg1139_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1139_out;
SharedReg1126_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1126_out;
SharedReg254_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg254_out;
SharedReg1155_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1155_out;
SharedReg1117_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1117_out;
SharedReg1118_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1118_out;
   MUX_Product18_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1119_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1125_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1117_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1118_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1131_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1121_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1123_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1141_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1139_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1126_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg254_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1155_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product18_1_impl_0_out);

   Delay1No370_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product18_1_impl_0_out,
                 Y => Delay1No370_out);

SharedReg854_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg854_out;
SharedReg1045_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1045_out;
SharedReg854_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg854_out;
SharedReg1081_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1081_out;
SharedReg158_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg158_out;
SharedReg672_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg672_out;
SharedReg674_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg674_out;
SharedReg1086_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1086_out;
SharedReg1115_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1115_out;
SharedReg746_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg746_out;
SharedReg337_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg337_out;
SharedReg374_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg374_out;
   MUX_Product18_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg854_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1045_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg337_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg374_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg854_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1081_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg158_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg672_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg674_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1086_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1115_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg746_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product18_1_impl_1_out);

   Delay1No371_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product18_1_impl_1_out,
                 Y => Delay1No371_out);

Delay1No372_out_to_Product18_2_impl_parent_implementedSystem_port_0_cast <= Delay1No372_out;
Delay1No373_out_to_Product18_2_impl_parent_implementedSystem_port_1_cast <= Delay1No373_out;
   Product18_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product18_2_impl_out,
                 X => Delay1No372_out_to_Product18_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No373_out_to_Product18_2_impl_parent_implementedSystem_port_1_cast);

SharedReg1117_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1117_out;
SharedReg1118_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1118_out;
SharedReg1119_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1125_out;
SharedReg1131_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1131_out;
SharedReg1121_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1121_out;
SharedReg1123_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1123_out;
SharedReg1141_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1141_out;
SharedReg1139_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1139_out;
SharedReg1126_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1126_out;
SharedReg260_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg260_out;
SharedReg1155_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1155_out;
   MUX_Product18_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1117_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1118_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg260_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1155_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1119_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1125_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1131_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1121_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1123_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1141_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1139_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1126_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product18_2_impl_0_out);

   Delay1No372_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product18_2_impl_0_out,
                 Y => Delay1No372_out);

SharedReg304_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg304_out;
SharedReg345_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg345_out;
SharedReg678_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg678_out;
SharedReg1015_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1015_out;
SharedReg678_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg678_out;
SharedReg1047_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1047_out;
SharedReg41_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg41_out;
SharedReg678_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg678_out;
SharedReg578_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg578_out;
SharedReg1052_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1052_out;
SharedReg1115_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1115_out;
SharedReg753_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg753_out;
   MUX_Product18_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg304_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg345_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1115_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg753_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg678_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1015_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg678_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1047_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg41_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg678_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg578_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1052_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product18_2_impl_1_out);

   Delay1No373_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product18_2_impl_1_out,
                 Y => Delay1No373_out);

Delay1No374_out_to_Product18_3_impl_parent_implementedSystem_port_0_cast <= Delay1No374_out;
Delay1No375_out_to_Product18_3_impl_parent_implementedSystem_port_1_cast <= Delay1No375_out;
   Product18_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product18_3_impl_out,
                 X => Delay1No374_out_to_Product18_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No375_out_to_Product18_3_impl_parent_implementedSystem_port_1_cast);

SharedReg1155_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1155_out;
SharedReg1117_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1117_out;
SharedReg1118_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1118_out;
SharedReg1119_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1125_out;
SharedReg1131_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1131_out;
SharedReg1121_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1121_out;
SharedReg1123_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1123_out;
SharedReg1141_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1141_out;
SharedReg1139_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1139_out;
SharedReg1126_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1126_out;
SharedReg266_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg266_out;
   MUX_Product18_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1155_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1117_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1126_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg266_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1118_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1119_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1125_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1131_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1121_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1123_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1141_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1139_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product18_3_impl_0_out);

   Delay1No374_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product18_3_impl_0_out,
                 Y => Delay1No374_out);

SharedReg758_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg758_out;
SharedReg352_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg352_out;
SharedReg193_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg193_out;
SharedReg683_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg683_out;
SharedReg1056_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1056_out;
SharedReg683_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg683_out;
SharedReg790_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg790_out;
SharedReg198_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg198_out;
SharedReg861_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg861_out;
SharedReg685_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg685_out;
SharedReg1058_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1058_out;
SharedReg1115_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1115_out;
   MUX_Product18_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg758_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg352_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1058_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1115_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg193_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg683_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1056_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg683_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg790_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg198_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg861_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg685_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product18_3_impl_1_out);

   Delay1No375_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product18_3_impl_1_out,
                 Y => Delay1No375_out);

Delay1No376_out_to_Product18_4_impl_parent_implementedSystem_port_0_cast <= Delay1No376_out;
Delay1No377_out_to_Product18_4_impl_parent_implementedSystem_port_1_cast <= Delay1No377_out;
   Product18_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product18_4_impl_out,
                 X => Delay1No376_out_to_Product18_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No377_out_to_Product18_4_impl_parent_implementedSystem_port_1_cast);

SharedReg1126_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1126_out;
SharedReg272_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg272_out;
SharedReg1155_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1155_out;
SharedReg1117_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1117_out;
SharedReg1118_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1118_out;
SharedReg1119_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1125_out;
SharedReg1131_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1131_out;
SharedReg1121_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1121_out;
SharedReg1123_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1123_out;
SharedReg1141_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1141_out;
SharedReg1139_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1139_out;
   MUX_Product18_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1126_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg272_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1141_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1139_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1155_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1117_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1118_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1119_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1125_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1131_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1121_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1123_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product18_4_impl_0_out);

   Delay1No376_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product18_4_impl_0_out,
                 Y => Delay1No376_out);

SharedReg1025_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1025_out;
SharedReg1115_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1115_out;
SharedReg764_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg764_out;
SharedReg310_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg310_out;
SharedReg281_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg281_out;
SharedReg584_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg584_out;
SharedReg995_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg995_out;
SharedReg689_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg689_out;
SharedReg764_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg764_out;
SharedReg48_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg48_out;
SharedReg689_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg689_out;
SharedReg691_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg691_out;
   MUX_Product18_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1025_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1115_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg689_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg691_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg764_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg310_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg281_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg584_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg995_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg689_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg764_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg48_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product18_4_impl_1_out);

   Delay1No377_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product18_4_impl_1_out,
                 Y => Delay1No377_out);

Delay1No378_out_to_Product18_5_impl_parent_implementedSystem_port_0_cast <= Delay1No378_out;
Delay1No379_out_to_Product18_5_impl_parent_implementedSystem_port_1_cast <= Delay1No379_out;
   Product18_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product18_5_impl_out,
                 X => Delay1No378_out_to_Product18_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No379_out_to_Product18_5_impl_parent_implementedSystem_port_1_cast);

SharedReg1141_out_to_MUX_Product18_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1141_out;
SharedReg1139_out_to_MUX_Product18_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1139_out;
SharedReg1126_out_to_MUX_Product18_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1126_out;
SharedReg212_out_to_MUX_Product18_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg212_out;
SharedReg1155_out_to_MUX_Product18_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1155_out;
SharedReg1117_out_to_MUX_Product18_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1117_out;
SharedReg1118_out_to_MUX_Product18_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1118_out;
SharedReg1119_out_to_MUX_Product18_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product18_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1125_out;
SharedReg1131_out_to_MUX_Product18_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1131_out;
SharedReg1121_out_to_MUX_Product18_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1121_out;
SharedReg1123_out_to_MUX_Product18_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1123_out;
   MUX_Product18_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1141_out_to_MUX_Product18_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1139_out_to_MUX_Product18_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1121_out_to_MUX_Product18_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1123_out_to_MUX_Product18_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1126_out_to_MUX_Product18_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg212_out_to_MUX_Product18_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1155_out_to_MUX_Product18_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1117_out_to_MUX_Product18_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1118_out_to_MUX_Product18_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1119_out_to_MUX_Product18_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1125_out_to_MUX_Product18_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1131_out_to_MUX_Product18_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product18_5_impl_0_out);

   Delay1No378_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product18_5_impl_0_out,
                 Y => Delay1No378_out);

SharedReg694_out_to_MUX_Product18_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg694_out;
SharedReg696_out_to_MUX_Product18_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg696_out;
SharedReg1063_out_to_MUX_Product18_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1063_out;
SharedReg1115_out_to_MUX_Product18_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1115_out;
SharedReg770_out_to_MUX_Product18_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg770_out;
SharedReg288_out_to_MUX_Product18_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg288_out;
SharedReg293_out_to_MUX_Product18_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg293_out;
SharedReg694_out_to_MUX_Product18_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg694_out;
SharedReg1000_out_to_MUX_Product18_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1000_out;
SharedReg868_out_to_MUX_Product18_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg868_out;
SharedReg770_out_to_MUX_Product18_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg770_out;
SharedReg118_out_to_MUX_Product18_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg118_out;
   MUX_Product18_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg694_out_to_MUX_Product18_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg696_out_to_MUX_Product18_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg770_out_to_MUX_Product18_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg118_out_to_MUX_Product18_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1063_out_to_MUX_Product18_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1115_out_to_MUX_Product18_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg770_out_to_MUX_Product18_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg288_out_to_MUX_Product18_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg293_out_to_MUX_Product18_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg694_out_to_MUX_Product18_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1000_out_to_MUX_Product18_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg868_out_to_MUX_Product18_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product18_5_impl_1_out);

   Delay1No379_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product18_5_impl_1_out,
                 Y => Delay1No379_out);

Delay1No380_out_to_Product18_6_impl_parent_implementedSystem_port_0_cast <= Delay1No380_out;
Delay1No381_out_to_Product18_6_impl_parent_implementedSystem_port_1_cast <= Delay1No381_out;
   Product18_6_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product18_6_impl_out,
                 X => Delay1No380_out_to_Product18_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No381_out_to_Product18_6_impl_parent_implementedSystem_port_1_cast);

SharedReg1123_out_to_MUX_Product18_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1123_out;
SharedReg1141_out_to_MUX_Product18_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1141_out;
SharedReg1139_out_to_MUX_Product18_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1139_out;
SharedReg1126_out_to_MUX_Product18_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1126_out;
SharedReg218_out_to_MUX_Product18_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg218_out;
SharedReg1155_out_to_MUX_Product18_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1155_out;
SharedReg1117_out_to_MUX_Product18_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1117_out;
SharedReg1118_out_to_MUX_Product18_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1118_out;
SharedReg1119_out_to_MUX_Product18_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product18_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1125_out;
SharedReg1131_out_to_MUX_Product18_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1131_out;
SharedReg1121_out_to_MUX_Product18_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1121_out;
   MUX_Product18_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1123_out_to_MUX_Product18_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1141_out_to_MUX_Product18_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1131_out_to_MUX_Product18_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1121_out_to_MUX_Product18_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1139_out_to_MUX_Product18_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1126_out_to_MUX_Product18_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg218_out_to_MUX_Product18_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1155_out_to_MUX_Product18_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1117_out_to_MUX_Product18_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1118_out_to_MUX_Product18_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1119_out_to_MUX_Product18_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1125_out_to_MUX_Product18_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product18_6_impl_0_out);

   Delay1No380_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product18_6_impl_0_out,
                 Y => Delay1No380_out);

SharedReg60_out_to_MUX_Product18_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg60_out;
SharedReg1001_out_to_MUX_Product18_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1001_out;
SharedReg1003_out_to_MUX_Product18_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1003_out;
SharedReg1093_out_to_MUX_Product18_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1093_out;
SharedReg1115_out_to_MUX_Product18_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1115_out;
SharedReg1088_out_to_MUX_Product18_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1088_out;
SharedReg322_out_to_MUX_Product18_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg322_out;
SharedReg358_out_to_MUX_Product18_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg358_out;
SharedReg1001_out_to_MUX_Product18_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1001_out;
SharedReg1078_out_to_MUX_Product18_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1078_out;
SharedReg1001_out_to_MUX_Product18_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1001_out;
SharedReg1101_out_to_MUX_Product18_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1101_out;
   MUX_Product18_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg60_out_to_MUX_Product18_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1001_out_to_MUX_Product18_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1001_out_to_MUX_Product18_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1101_out_to_MUX_Product18_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1003_out_to_MUX_Product18_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1093_out_to_MUX_Product18_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1115_out_to_MUX_Product18_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1088_out_to_MUX_Product18_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg322_out_to_MUX_Product18_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg358_out_to_MUX_Product18_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1001_out_to_MUX_Product18_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1078_out_to_MUX_Product18_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product18_6_impl_1_out);

   Delay1No381_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product18_6_impl_1_out,
                 Y => Delay1No381_out);

Delay1No382_out_to_Product28_0_impl_parent_implementedSystem_port_0_cast <= Delay1No382_out;
Delay1No383_out_to_Product28_0_impl_parent_implementedSystem_port_1_cast <= Delay1No383_out;
   Product28_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product28_0_impl_out,
                 X => Delay1No382_out_to_Product28_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No383_out_to_Product28_0_impl_parent_implementedSystem_port_1_cast);

SharedReg1004_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1004_out;
SharedReg1038_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1038_out;
SharedReg127_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg127_out;
SharedReg981_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg981_out;
SharedReg983_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg983_out;
SharedReg1098_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1098_out;
SharedReg1103_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1103_out;
SharedReg1157_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1157_out;
SharedReg1105_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1105_out;
SharedReg203_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg203_out;
SharedReg1004_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1004_out;
SharedReg1097_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1097_out;
   MUX_Product28_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1004_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1038_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1004_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1097_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg127_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg981_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg983_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1098_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1103_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1157_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1105_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg203_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product28_0_impl_0_out);

   Delay1No382_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_0_impl_0_out,
                 Y => Delay1No382_out);

SharedReg1131_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1131_out;
SharedReg1121_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1121_out;
SharedReg1123_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1123_out;
SharedReg1141_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1141_out;
SharedReg1139_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1139_out;
SharedReg1126_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1126_out;
SharedReg363_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg363_out;
SharedReg775_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg775_out;
SharedReg128_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg128_out;
SharedReg1118_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1118_out;
SharedReg1119_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1125_out;
   MUX_Product28_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1131_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1121_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1119_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1125_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1123_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1141_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1139_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1126_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg363_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg775_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg128_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1118_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product28_0_impl_1_out);

   Delay1No383_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_0_impl_1_out,
                 Y => Delay1No383_out);

Delay1No384_out_to_Product28_1_impl_parent_implementedSystem_port_0_cast <= Delay1No384_out;
Delay1No385_out_to_Product28_1_impl_parent_implementedSystem_port_1_cast <= Delay1No385_out;
   Product28_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product28_1_impl_out,
                 X => Delay1No384_out_to_Product28_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No385_out_to_Product28_1_impl_parent_implementedSystem_port_1_cast);

SharedReg984_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg984_out;
SharedReg1084_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1084_out;
SharedReg984_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg984_out;
SharedReg1008_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1008_out;
SharedReg100_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg100_out;
SharedReg854_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg854_out;
SharedReg856_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg856_out;
SharedReg1085_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1085_out;
SharedReg1103_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1103_out;
SharedReg1157_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1157_out;
SharedReg1105_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1105_out;
SharedReg236_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg236_out;
   MUX_Product28_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg984_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1084_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1105_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg236_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg984_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1008_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg100_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg854_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg856_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1085_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1103_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1157_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product28_1_impl_0_out);

   Delay1No384_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_1_impl_0_out,
                 Y => Delay1No384_out);

SharedReg1119_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1125_out;
SharedReg1131_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1131_out;
SharedReg1121_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1121_out;
SharedReg1123_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1123_out;
SharedReg1141_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1141_out;
SharedReg1139_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1139_out;
SharedReg1126_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1126_out;
SharedReg164_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg164_out;
SharedReg746_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg746_out;
SharedReg131_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg131_out;
SharedReg1118_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1118_out;
   MUX_Product28_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1119_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1125_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg131_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1118_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1131_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1121_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1123_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1141_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1139_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1126_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg164_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg746_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product28_1_impl_1_out);

   Delay1No385_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_1_impl_1_out,
                 Y => Delay1No385_out);

Delay1No386_out_to_Product28_2_impl_parent_implementedSystem_port_0_cast <= Delay1No386_out;
Delay1No387_out_to_Product28_2_impl_parent_implementedSystem_port_1_cast <= Delay1No387_out;
   Product28_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product28_2_impl_out,
                 X => Delay1No386_out_to_Product28_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No387_out_to_Product28_2_impl_parent_implementedSystem_port_1_cast);

SharedReg1105_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1105_out;
SharedReg241_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg241_out;
SharedReg858_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg858_out;
SharedReg1050_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1050_out;
SharedReg858_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg858_out;
SharedReg987_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg987_out;
SharedReg134_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg134_out;
SharedReg858_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg858_out;
SharedReg680_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg680_out;
SharedReg1051_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1051_out;
SharedReg1103_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1103_out;
SharedReg1157_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1157_out;
   MUX_Product28_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1105_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg241_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1103_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1157_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg858_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1050_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg858_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg987_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg134_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg858_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg680_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1051_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product28_2_impl_0_out);

   Delay1No386_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_2_impl_0_out,
                 Y => Delay1No386_out);

SharedReg135_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg135_out;
SharedReg1118_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1118_out;
SharedReg1119_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1125_out;
SharedReg1131_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1131_out;
SharedReg1121_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1121_out;
SharedReg1123_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1123_out;
SharedReg1141_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1141_out;
SharedReg1139_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1139_out;
SharedReg1126_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1126_out;
SharedReg170_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg170_out;
SharedReg753_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg753_out;
   MUX_Product28_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg135_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1118_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg170_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg753_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1119_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1125_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1131_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1121_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1123_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1141_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1139_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1126_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product28_2_impl_1_out);

   Delay1No387_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_2_impl_1_out,
                 Y => Delay1No387_out);

Delay1No388_out_to_Product28_3_impl_parent_implementedSystem_port_0_cast <= Delay1No388_out;
Delay1No389_out_to_Product28_3_impl_parent_implementedSystem_port_1_cast <= Delay1No389_out;
   Product28_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product28_3_impl_out,
                 X => Delay1No388_out_to_Product28_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No389_out_to_Product28_3_impl_parent_implementedSystem_port_1_cast);

SharedReg1157_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1157_out;
SharedReg1105_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1105_out;
SharedReg141_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg141_out;
SharedReg861_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg861_out;
SharedReg793_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg793_out;
SharedReg861_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg861_out;
SharedReg991_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg991_out;
SharedReg110_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg110_out;
SharedReg990_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg990_out;
SharedReg863_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg863_out;
SharedReg1057_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1057_out;
SharedReg1103_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1103_out;
   MUX_Product28_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1157_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1105_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1057_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1103_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg141_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg861_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg793_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg861_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg991_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg110_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg990_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg863_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product28_3_impl_0_out);

   Delay1No388_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_3_impl_0_out,
                 Y => Delay1No388_out);

SharedReg758_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg758_out;
SharedReg111_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg111_out;
SharedReg1118_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1118_out;
SharedReg1119_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1125_out;
SharedReg1131_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1131_out;
SharedReg1121_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1121_out;
SharedReg1123_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1123_out;
SharedReg1141_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1141_out;
SharedReg1139_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1139_out;
SharedReg1126_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1126_out;
SharedReg175_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg175_out;
   MUX_Product28_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg758_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg111_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1126_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg175_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1118_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1119_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1125_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1131_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1121_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1123_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1141_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1139_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product28_3_impl_1_out);

   Delay1No389_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_3_impl_1_out,
                 Y => Delay1No389_out);

Delay1No390_out_to_Product28_4_impl_parent_implementedSystem_port_0_cast <= Delay1No390_out;
Delay1No391_out_to_Product28_4_impl_parent_implementedSystem_port_1_cast <= Delay1No391_out;
   Product28_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product28_4_impl_out,
                 X => Delay1No390_out_to_Product28_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No391_out_to_Product28_4_impl_parent_implementedSystem_port_1_cast);

SharedReg799_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg799_out;
SharedReg1103_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1103_out;
SharedReg1157_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1157_out;
SharedReg1105_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1105_out;
SharedReg147_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg147_out;
SharedReg689_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg689_out;
SharedReg1024_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1024_out;
SharedReg865_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg865_out;
SharedReg994_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg994_out;
SharedReg145_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg145_out;
SharedReg865_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg865_out;
SharedReg867_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg867_out;
   MUX_Product28_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg799_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1103_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg865_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg867_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1157_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1105_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg147_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg689_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1024_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg865_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg994_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg145_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product28_4_impl_0_out);

   Delay1No390_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_4_impl_0_out,
                 Y => Delay1No390_out);

SharedReg1126_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1126_out;
SharedReg52_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg52_out;
SharedReg764_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg764_out;
SharedReg115_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg115_out;
SharedReg1118_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1118_out;
SharedReg1119_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1125_out;
SharedReg1131_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1131_out;
SharedReg1121_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1121_out;
SharedReg1123_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1123_out;
SharedReg1141_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1141_out;
SharedReg1139_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1139_out;
   MUX_Product28_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1126_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg52_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1141_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1139_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg764_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg115_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1118_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1119_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1125_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1131_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1121_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1123_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product28_4_impl_1_out);

   Delay1No391_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_4_impl_1_out,
                 Y => Delay1No391_out);

Delay1No392_out_to_Product28_5_impl_parent_implementedSystem_port_0_cast <= Delay1No392_out;
Delay1No393_out_to_Product28_5_impl_parent_implementedSystem_port_1_cast <= Delay1No393_out;
   Product28_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product28_5_impl_out,
                 X => Delay1No392_out_to_Product28_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No393_out_to_Product28_5_impl_parent_implementedSystem_port_1_cast);

SharedReg868_out_to_MUX_Product28_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg868_out;
SharedReg870_out_to_MUX_Product28_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg870_out;
SharedReg774_out_to_MUX_Product28_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg774_out;
SharedReg1103_out_to_MUX_Product28_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1103_out;
SharedReg1157_out_to_MUX_Product28_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1157_out;
SharedReg1105_out_to_MUX_Product28_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1105_out;
SharedReg184_out_to_MUX_Product28_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg184_out;
SharedReg868_out_to_MUX_Product28_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg868_out;
SharedReg1031_out_to_MUX_Product28_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1031_out;
SharedReg997_out_to_MUX_Product28_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg997_out;
SharedReg1029_out_to_MUX_Product28_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1029_out;
SharedReg212_out_to_MUX_Product28_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg212_out;
   MUX_Product28_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg868_out_to_MUX_Product28_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg870_out_to_MUX_Product28_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1029_out_to_MUX_Product28_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg212_out_to_MUX_Product28_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg774_out_to_MUX_Product28_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1103_out_to_MUX_Product28_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1157_out_to_MUX_Product28_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1105_out_to_MUX_Product28_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg184_out_to_MUX_Product28_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg868_out_to_MUX_Product28_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1031_out_to_MUX_Product28_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg997_out_to_MUX_Product28_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product28_5_impl_0_out);

   Delay1No392_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_5_impl_0_out,
                 Y => Delay1No392_out);

SharedReg1141_out_to_MUX_Product28_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1141_out;
SharedReg1139_out_to_MUX_Product28_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1139_out;
SharedReg1126_out_to_MUX_Product28_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1126_out;
SharedReg313_out_to_MUX_Product28_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg313_out;
SharedReg770_out_to_MUX_Product28_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg770_out;
SharedReg151_out_to_MUX_Product28_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg151_out;
SharedReg1118_out_to_MUX_Product28_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1118_out;
SharedReg1119_out_to_MUX_Product28_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product28_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1125_out;
SharedReg1131_out_to_MUX_Product28_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1131_out;
SharedReg1121_out_to_MUX_Product28_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1121_out;
SharedReg1123_out_to_MUX_Product28_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1123_out;
   MUX_Product28_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1141_out_to_MUX_Product28_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1139_out_to_MUX_Product28_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1121_out_to_MUX_Product28_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1123_out_to_MUX_Product28_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1126_out_to_MUX_Product28_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg313_out_to_MUX_Product28_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg770_out_to_MUX_Product28_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg151_out_to_MUX_Product28_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1118_out_to_MUX_Product28_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1119_out_to_MUX_Product28_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1125_out_to_MUX_Product28_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1131_out_to_MUX_Product28_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product28_5_impl_1_out);

   Delay1No393_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_5_impl_1_out,
                 Y => Delay1No393_out);

Delay1No394_out_to_Product28_6_impl_parent_implementedSystem_port_0_cast <= Delay1No394_out;
Delay1No395_out_to_Product28_6_impl_parent_implementedSystem_port_1_cast <= Delay1No395_out;
   Product28_6_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product28_6_impl_out,
                 X => Delay1No394_out_to_Product28_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No395_out_to_Product28_6_impl_parent_implementedSystem_port_1_cast);

SharedReg153_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg153_out;
SharedReg1033_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1033_out;
SharedReg1036_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1036_out;
SharedReg1092_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1092_out;
SharedReg1103_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1103_out;
SharedReg1157_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1157_out;
SharedReg1105_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1105_out;
SharedReg155_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg155_out;
SharedReg1033_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1033_out;
SharedReg1091_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1091_out;
SharedReg1033_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1033_out;
SharedReg1067_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1067_out;
   MUX_Product28_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg153_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1033_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1033_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1067_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1036_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1092_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1103_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1157_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1105_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg155_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1033_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1091_out_to_MUX_Product28_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product28_6_impl_0_out);

   Delay1No394_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_6_impl_0_out,
                 Y => Delay1No394_out);

SharedReg1123_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1123_out;
SharedReg1141_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1141_out;
SharedReg1139_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1139_out;
SharedReg1126_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1126_out;
SharedReg381_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg381_out;
SharedReg1088_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1088_out;
SharedReg124_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg124_out;
SharedReg1118_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1118_out;
SharedReg1119_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1119_out;
SharedReg1125_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1125_out;
SharedReg1131_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1131_out;
SharedReg1121_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1121_out;
   MUX_Product28_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1123_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1141_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1131_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1121_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1139_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1126_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg381_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1088_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg124_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1118_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1119_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1125_out_to_MUX_Product28_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product28_6_impl_1_out);

   Delay1No395_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_6_impl_1_out,
                 Y => Delay1No395_out);

Delay1No396_out_to_Subtract9_0_impl_parent_implementedSystem_port_0_cast <= Delay1No396_out;
Delay1No397_out_to_Subtract9_0_impl_parent_implementedSystem_port_1_cast <= Delay1No397_out;
   Subtract9_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract9_0_impl_out,
                 X => Delay1No396_out_to_Subtract9_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No397_out_to_Subtract9_0_impl_parent_implementedSystem_port_1_cast);

SharedReg886_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg886_out;
SharedReg3_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg3_out;
SharedReg940_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg940_out;
SharedReg646_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg646_out;
SharedReg883_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg883_out;
SharedReg883_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg883_out;
SharedReg251_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg251_out;
SharedReg564_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg564_out;
SharedReg434_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg434_out;
SharedReg666_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg666_out;
SharedReg850_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg850_out;
SharedReg800_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg800_out;
   MUX_Subtract9_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg886_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg3_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg850_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg800_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg940_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg646_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg883_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg883_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg251_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg564_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg434_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg666_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract9_0_impl_0_out);

   Delay1No396_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_0_impl_0_out,
                 Y => Delay1No396_out);

Delay4No266_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_1_cast <= Delay4No266_out;
SharedReg19_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg19_out;
SharedReg941_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg941_out;
SharedReg822_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg822_out;
SharedReg960_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg960_out;
SharedReg960_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg960_out;
SharedReg334_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg334_out;
SharedReg849_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg849_out;
SharedReg1037_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1037_out;
SharedReg982_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg982_out;
SharedReg849_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg849_out;
SharedReg604_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg604_out;
   MUX_Subtract9_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay4No266_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg19_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg849_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg604_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg941_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg822_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg960_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg960_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg334_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg849_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1037_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg982_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract9_0_impl_1_out);

   Delay1No397_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_0_impl_1_out,
                 Y => Delay1No397_out);

Delay1No398_out_to_Subtract9_1_impl_parent_implementedSystem_port_0_cast <= Delay1No398_out;
Delay1No399_out_to_Subtract9_1_impl_parent_implementedSystem_port_1_cast <= Delay1No399_out;
   Subtract9_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract9_1_impl_out,
                 X => Delay1No398_out_to_Subtract9_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No399_out_to_Subtract9_1_impl_parent_implementedSystem_port_1_cast);

SharedReg235_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg235_out;
SharedReg803_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg803_out;
SharedReg890_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg890_out;
SharedReg3_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg3_out;
SharedReg943_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg943_out;
SharedReg888_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg888_out;
SharedReg533_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg533_out;
SharedReg1007_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1007_out;
SharedReg1044_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1044_out;
SharedReg1084_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1084_out;
SharedReg338_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg338_out;
SharedReg130_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg130_out;
   MUX_Subtract9_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg235_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg803_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg338_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg130_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg890_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg3_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg943_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg888_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg533_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1007_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1044_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1084_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract9_1_impl_0_out);

   Delay1No398_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_1_impl_0_out,
                 Y => Delay1No398_out);

SharedReg372_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg372_out;
SharedReg607_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg607_out;
Delay4No267_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_3_cast <= Delay4No267_out;
SharedReg19_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg19_out;
SharedReg944_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg944_out;
SharedReg964_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg964_out;
SharedReg628_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg628_out;
SharedReg570_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg570_out;
SharedReg574_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg574_out;
SharedReg438_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg438_out;
SharedReg372_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg372_out;
SharedReg336_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg336_out;
   MUX_Subtract9_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg372_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg607_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg372_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg336_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => Delay4No267_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg19_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg944_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg964_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg628_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg570_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg574_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg438_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract9_1_impl_1_out);

   Delay1No399_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_1_impl_1_out,
                 Y => Delay1No399_out);

Delay1No400_out_to_Subtract9_2_impl_parent_implementedSystem_port_0_cast <= Delay1No400_out;
Delay1No401_out_to_Subtract9_2_impl_parent_implementedSystem_port_1_cast <= Delay1No401_out;
   Subtract9_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract9_2_impl_out,
                 X => Delay1No400_out_to_Subtract9_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No401_out_to_Subtract9_2_impl_parent_implementedSystem_port_1_cast);

SharedReg343_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg343_out;
SharedReg134_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg134_out;
SharedReg240_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg240_out;
SharedReg806_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg806_out;
SharedReg894_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg894_out;
SharedReg4_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg7_out;
SharedReg611_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg611_out;
SharedReg652_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg652_out;
SharedReg171_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg171_out;
SharedReg344_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg344_out;
SharedReg200_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg200_out;
   MUX_Subtract9_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg343_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg134_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg344_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg200_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg240_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg806_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg894_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg4_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg7_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg611_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg652_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg171_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract9_2_impl_0_out);

   Delay1No400_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_2_impl_0_out,
                 Y => Delay1No400_out);

SharedReg170_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg170_out;
SharedReg303_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg303_out;
SharedReg342_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg342_out;
SharedReg610_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg610_out;
Delay4No268_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_5_cast <= Delay4No268_out;
SharedReg20_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg20_out;
SharedReg23_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg23_out;
SharedReg894_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg894_out;
SharedReg830_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg830_out;
SharedReg342_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg342_out;
SharedReg348_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg348_out;
SharedReg302_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg302_out;
   MUX_Subtract9_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg170_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg303_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg348_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg302_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg342_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg610_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay4No268_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg20_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg23_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg894_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg830_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg342_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract9_2_impl_1_out);

   Delay1No401_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_2_impl_1_out,
                 Y => Delay1No401_out);

Delay1No402_out_to_Subtract9_3_impl_parent_implementedSystem_port_0_cast <= Delay1No402_out;
Delay1No403_out_to_Subtract9_3_impl_parent_implementedSystem_port_1_cast <= Delay1No403_out;
   Subtract9_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract9_3_impl_out,
                 X => Delay1No402_out_to_Subtract9_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No403_out_to_Subtract9_3_impl_parent_implementedSystem_port_1_cast);

SharedReg178_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg178_out;
SharedReg194_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg194_out;
SharedReg110_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg110_out;
SharedReg581_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg581_out;
SharedReg809_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg809_out;
SharedReg898_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg898_out;
SharedReg3_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg3_out;
SharedReg7_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg7_out;
SharedReg896_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg896_out;
SharedReg655_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg655_out;
SharedReg192_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg192_out;
SharedReg352_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg352_out;
   MUX_Subtract9_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg178_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg194_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg192_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg352_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg110_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg581_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg809_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg898_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg3_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg7_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg896_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg655_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract9_3_impl_0_out);

   Delay1No402_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_3_impl_0_out,
                 Y => Delay1No402_out);

SharedReg266_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg266_out;
SharedReg191_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg191_out;
SharedReg351_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg351_out;
SharedReg580_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg580_out;
SharedReg613_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg613_out;
Delay4No269_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_6_cast <= Delay4No269_out;
SharedReg19_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg19_out;
SharedReg23_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg23_out;
SharedReg970_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg970_out;
SharedReg834_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg834_out;
SharedReg350_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg350_out;
SharedReg354_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg354_out;
   MUX_Subtract9_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg266_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg191_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg350_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg354_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg351_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg580_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg613_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay4No269_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg19_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg23_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg970_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg834_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract9_3_impl_1_out);

   Delay1No403_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_3_impl_1_out,
                 Y => Delay1No403_out);

Delay1No404_out_to_Subtract9_4_impl_parent_implementedSystem_port_0_cast <= Delay1No404_out;
Delay1No405_out_to_Subtract9_4_impl_parent_implementedSystem_port_1_cast <= Delay1No405_out;
   Subtract9_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract9_4_impl_out,
                 X => Delay1No404_out_to_Subtract9_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No405_out_to_Subtract9_4_impl_parent_implementedSystem_port_1_cast);

SharedReg705_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg705_out;
SharedReg280_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg280_out;
SharedReg89_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg89_out;
SharedReg282_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg282_out;
SharedReg114_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg114_out;
SharedReg146_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg146_out;
SharedReg812_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg812_out;
SharedReg56_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg56_out;
SharedReg4_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg4_out;
SharedReg8_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg8_out;
SharedReg901_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg901_out;
SharedReg408_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg408_out;
   MUX_Subtract9_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg705_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg280_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg901_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg408_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg89_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg282_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg114_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg146_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg812_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg56_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg4_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg8_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract9_4_impl_0_out);

   Delay1No404_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_4_impl_0_out,
                 Y => Delay1No404_out);

SharedReg866_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg866_out;
SharedReg285_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg285_out;
SharedReg272_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg272_out;
SharedReg308_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg308_out;
SharedReg273_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg273_out;
SharedReg308_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg308_out;
SharedReg616_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg616_out;
SharedReg59_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg59_out;
SharedReg20_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg20_out;
SharedReg24_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg24_out;
Delay5No46_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_11_cast <= Delay5No46_out;
SharedReg518_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg518_out;
   MUX_Subtract9_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg866_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg285_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay5No46_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg518_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg272_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg308_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg273_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg308_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg616_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg59_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg20_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg24_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract9_4_impl_1_out);

   Delay1No405_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_4_impl_1_out,
                 Y => Delay1No405_out);

Delay1No406_out_to_Subtract9_5_impl_parent_implementedSystem_port_0_cast <= Delay1No406_out;
Delay1No407_out_to_Subtract9_5_impl_parent_implementedSystem_port_1_cast <= Delay1No407_out;
   Subtract9_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract9_5_impl_out,
                 X => Delay1No406_out_to_Subtract9_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No407_out_to_Subtract9_5_impl_parent_implementedSystem_port_1_cast);

SharedReg905_out_to_MUX_Subtract9_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg905_out;
SharedReg661_out_to_MUX_Subtract9_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg661_out;
SharedReg225_out_to_MUX_Subtract9_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg225_out;
SharedReg1061_out_to_MUX_Subtract9_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1061_out;
SharedReg773_out_to_MUX_Subtract9_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg773_out;
SharedReg316_out_to_MUX_Subtract9_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg316_out;
SharedReg464_out_to_MUX_Subtract9_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg464_out;
SharedReg213_out_to_MUX_Subtract9_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg213_out;
SharedReg815_out_to_MUX_Subtract9_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg815_out;
SharedReg228_out_to_MUX_Subtract9_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg228_out;
SharedReg5_out_to_MUX_Subtract9_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg5_out;
SharedReg8_out_to_MUX_Subtract9_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg8_out;
   MUX_Subtract9_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg905_out_to_MUX_Subtract9_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg661_out_to_MUX_Subtract9_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg5_out_to_MUX_Subtract9_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg8_out_to_MUX_Subtract9_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg225_out_to_MUX_Subtract9_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1061_out_to_MUX_Subtract9_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg773_out_to_MUX_Subtract9_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg316_out_to_MUX_Subtract9_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg464_out_to_MUX_Subtract9_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg213_out_to_MUX_Subtract9_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg815_out_to_MUX_Subtract9_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg228_out_to_MUX_Subtract9_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract9_5_impl_0_out);

   Delay1No406_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_5_impl_0_out,
                 Y => Delay1No406_out);

Delay5No47_out_to_MUX_Subtract9_5_impl_1_parent_implementedSystem_port_1_cast <= Delay5No47_out;
SharedReg842_out_to_MUX_Subtract9_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg842_out;
SharedReg290_out_to_MUX_Subtract9_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg290_out;
SharedReg593_out_to_MUX_Subtract9_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg593_out;
SharedReg764_out_to_MUX_Subtract9_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg764_out;
SharedReg290_out_to_MUX_Subtract9_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg290_out;
SharedReg590_out_to_MUX_Subtract9_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg590_out;
SharedReg313_out_to_MUX_Subtract9_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg313_out;
SharedReg619_out_to_MUX_Subtract9_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg619_out;
SharedReg233_out_to_MUX_Subtract9_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg233_out;
SharedReg21_out_to_MUX_Subtract9_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg21_out;
SharedReg24_out_to_MUX_Subtract9_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg24_out;
   MUX_Subtract9_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay5No47_out_to_MUX_Subtract9_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg842_out_to_MUX_Subtract9_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg21_out_to_MUX_Subtract9_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg24_out_to_MUX_Subtract9_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg290_out_to_MUX_Subtract9_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg593_out_to_MUX_Subtract9_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg764_out_to_MUX_Subtract9_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg290_out_to_MUX_Subtract9_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg590_out_to_MUX_Subtract9_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg313_out_to_MUX_Subtract9_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg619_out_to_MUX_Subtract9_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg233_out_to_MUX_Subtract9_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract9_5_impl_1_out);

   Delay1No407_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_5_impl_1_out,
                 Y => Delay1No407_out);

Delay1No408_out_to_Subtract9_6_impl_parent_implementedSystem_port_0_cast <= Delay1No408_out;
Delay1No409_out_to_Subtract9_6_impl_parent_implementedSystem_port_1_cast <= Delay1No409_out;
   Subtract9_6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract9_6_impl_out,
                 X => Delay1No408_out_to_Subtract9_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No409_out_to_Subtract9_6_impl_parent_implementedSystem_port_1_cast);

SharedReg7_out_to_MUX_Subtract9_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg7_out;
SharedReg664_out_to_MUX_Subtract9_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg664_out;
SharedReg548_out_to_MUX_Subtract9_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg548_out;
SharedReg907_out_to_MUX_Subtract9_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg907_out;
SharedReg220_out_to_MUX_Subtract9_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg220_out;
SharedReg473_out_to_MUX_Subtract9_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg473_out;
SharedReg908_out_to_MUX_Subtract9_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg908_out;
SharedReg595_out_to_MUX_Subtract9_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg595_out;
SharedReg92_out_to_MUX_Subtract9_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg92_out;
SharedReg818_out_to_MUX_Subtract9_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg818_out;
SharedReg910_out_to_MUX_Subtract9_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg910_out;
SharedReg3_out_to_MUX_Subtract9_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg3_out;
   MUX_Subtract9_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg7_out_to_MUX_Subtract9_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg664_out_to_MUX_Subtract9_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg910_out_to_MUX_Subtract9_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg3_out_to_MUX_Subtract9_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg548_out_to_MUX_Subtract9_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg907_out_to_MUX_Subtract9_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg220_out_to_MUX_Subtract9_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg473_out_to_MUX_Subtract9_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg908_out_to_MUX_Subtract9_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg595_out_to_MUX_Subtract9_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg92_out_to_MUX_Subtract9_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg818_out_to_MUX_Subtract9_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract9_6_impl_0_out);

   Delay1No408_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_6_impl_0_out,
                 Y => Delay1No408_out);

SharedReg23_out_to_MUX_Subtract9_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg23_out;
SharedReg846_out_to_MUX_Subtract9_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg846_out;
SharedReg643_out_to_MUX_Subtract9_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg643_out;
SharedReg978_out_to_MUX_Subtract9_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg978_out;
SharedReg362_out_to_MUX_Subtract9_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg362_out;
SharedReg699_out_to_MUX_Subtract9_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg699_out;
SharedReg979_out_to_MUX_Subtract9_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg979_out;
SharedReg1002_out_to_MUX_Subtract9_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1002_out;
SharedReg320_out_to_MUX_Subtract9_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg320_out;
SharedReg622_out_to_MUX_Subtract9_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg622_out;
Delay4No272_out_to_MUX_Subtract9_6_impl_1_parent_implementedSystem_port_11_cast <= Delay4No272_out;
SharedReg19_out_to_MUX_Subtract9_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg19_out;
   MUX_Subtract9_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg23_out_to_MUX_Subtract9_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg846_out_to_MUX_Subtract9_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay4No272_out_to_MUX_Subtract9_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg19_out_to_MUX_Subtract9_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg643_out_to_MUX_Subtract9_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg978_out_to_MUX_Subtract9_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg362_out_to_MUX_Subtract9_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg699_out_to_MUX_Subtract9_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg979_out_to_MUX_Subtract9_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1002_out_to_MUX_Subtract9_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg320_out_to_MUX_Subtract9_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg622_out_to_MUX_Subtract9_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract9_6_impl_1_out);

   Delay1No409_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_6_impl_1_out,
                 Y => Delay1No409_out);

Delay1No410_out_to_Subtract10_3_impl_parent_implementedSystem_port_0_cast <= Delay1No410_out;
Delay1No411_out_to_Subtract10_3_impl_parent_implementedSystem_port_1_cast <= Delay1No411_out;
   Subtract10_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract10_3_impl_out,
                 X => Delay1No410_out_to_Subtract10_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No411_out_to_Subtract10_3_impl_parent_implementedSystem_port_1_cast);

SharedReg404_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg404_out;
SharedReg302_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg302_out;
SharedReg171_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg171_out;
SharedReg946_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg946_out;
SharedReg173_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg173_out;
SharedReg13_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg13_out;
SharedReg12_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg12_out;
SharedReg263_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg263_out;
SharedReg579_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg579_out;
SharedReg404_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg404_out;
SharedReg404_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg404_out;
SharedReg404_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg404_out;
   MUX_Subtract10_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg404_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg302_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg404_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg404_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg171_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg946_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg173_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg13_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg12_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg263_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg579_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg404_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract10_3_impl_0_out);

   Delay1No410_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract10_3_impl_0_out,
                 Y => Delay1No410_out);

SharedReg513_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg513_out;
SharedReg264_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg264_out;
SharedReg347_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg347_out;
SharedReg966_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg966_out;
SharedReg265_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg265_out;
SharedReg29_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg29_out;
SharedReg28_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg28_out;
SharedReg304_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg304_out;
SharedReg748_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg748_out;
SharedReg513_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg513_out;
SharedReg513_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg513_out;
SharedReg513_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg513_out;
   MUX_Subtract10_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg513_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg264_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg513_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg513_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg347_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg966_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg265_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg29_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg28_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg304_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg748_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg513_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract10_3_impl_1_out);

   Delay1No411_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract10_3_impl_1_out,
                 Y => Delay1No411_out);

Delay1No412_out_to_Product50_0_impl_parent_implementedSystem_port_0_cast <= Delay1No412_out;
Delay1No413_out_to_Product50_0_impl_parent_implementedSystem_port_1_cast <= Delay1No413_out;
   Product50_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product50_0_impl_out,
                 X => Delay1No412_out_to_Product50_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No413_out_to_Product50_0_impl_parent_implementedSystem_port_1_cast);

SharedReg1129_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1129_out;
SharedReg1149_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1149_out;
SharedReg1136_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1136_out;
SharedReg1137_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1137_out;
SharedReg1135_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1135_out;
SharedReg1114_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1114_out;
SharedReg1115_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1115_out;
SharedReg364_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg364_out;
SharedReg128_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg128_out;
SharedReg1106_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1106_out;
SharedReg1148_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1148_out;
SharedReg1113_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1113_out;
   MUX_Product50_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1129_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1149_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1148_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1113_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1136_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1137_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1135_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1114_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1115_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg364_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg128_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1106_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product50_0_impl_0_out);

   Delay1No412_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product50_0_impl_0_out,
                 Y => Delay1No412_out);

SharedReg1070_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1070_out;
SharedReg850_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg850_out;
SharedReg849_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg849_out;
SharedReg564_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg564_out;
SharedReg1040_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1040_out;
SharedReg1100_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1100_out;
SharedReg430_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg430_out;
SharedReg1116_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1116_out;
SharedReg1117_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1117_out;
SharedReg34_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg34_out;
SharedReg1037_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1037_out;
SharedReg777_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg777_out;
   MUX_Product50_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1070_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg850_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1037_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg777_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg849_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg564_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1040_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1100_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg430_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1116_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1117_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg34_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product50_0_impl_1_out);

   Delay1No413_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product50_0_impl_1_out,
                 Y => Delay1No413_out);

Delay1No414_out_to_Product50_1_impl_parent_implementedSystem_port_0_cast <= Delay1No414_out;
Delay1No415_out_to_Product50_1_impl_parent_implementedSystem_port_1_cast <= Delay1No415_out;
   Product50_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product50_1_impl_out,
                 X => Delay1No414_out_to_Product50_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No415_out_to_Product50_1_impl_parent_implementedSystem_port_1_cast);

SharedReg1148_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1148_out;
SharedReg1113_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1113_out;
SharedReg1129_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1129_out;
SharedReg1149_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1149_out;
SharedReg1136_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1136_out;
SharedReg1137_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1137_out;
SharedReg1135_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1135_out;
SharedReg1114_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1114_out;
SharedReg1115_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1115_out;
SharedReg165_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg165_out;
SharedReg131_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg131_out;
SharedReg1106_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1106_out;
   MUX_Product50_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1148_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1113_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg131_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1106_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1129_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1149_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1136_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1137_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1135_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1114_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1115_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg165_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product50_1_impl_0_out);

   Delay1No414_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product50_1_impl_0_out,
                 Y => Delay1No414_out);

SharedReg1007_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1007_out;
SharedReg785_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg785_out;
SharedReg1042_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1042_out;
SharedReg673_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg673_out;
SharedReg672_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg672_out;
SharedReg438_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg438_out;
SharedReg1010_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1010_out;
SharedReg1087_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1087_out;
SharedReg438_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg438_out;
SharedReg1116_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1116_out;
SharedReg1117_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1117_out;
SharedReg39_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg39_out;
   MUX_Product50_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1007_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg785_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1117_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg39_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1042_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg673_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg672_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg438_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1010_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1087_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg438_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1116_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product50_1_impl_1_out);

   Delay1No415_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product50_1_impl_1_out,
                 Y => Delay1No415_out);

Delay1No416_out_to_Product50_2_impl_parent_implementedSystem_port_0_cast <= Delay1No416_out;
Delay1No417_out_to_Product50_2_impl_parent_implementedSystem_port_1_cast <= Delay1No417_out;
   Product50_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product50_2_impl_out,
                 X => Delay1No416_out_to_Product50_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No417_out_to_Product50_2_impl_parent_implementedSystem_port_1_cast);

SharedReg135_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg135_out;
SharedReg1106_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1106_out;
SharedReg1148_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1148_out;
SharedReg1113_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1113_out;
SharedReg1129_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1129_out;
SharedReg1149_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1149_out;
SharedReg1136_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1136_out;
SharedReg1137_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1137_out;
SharedReg1135_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1135_out;
SharedReg1114_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1114_out;
SharedReg1115_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1115_out;
SharedReg171_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg171_out;
   MUX_Product50_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg135_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1106_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1115_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg171_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1148_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1113_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1129_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1149_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1136_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1137_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1135_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1114_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product50_2_impl_0_out);

   Delay1No416_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product50_2_impl_0_out,
                 Y => Delay1No416_out);

SharedReg1117_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1117_out;
SharedReg42_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg42_out;
SharedReg986_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg986_out;
SharedReg878_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg878_out;
SharedReg1012_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1012_out;
SharedReg577_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg577_out;
SharedReg678_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg678_out;
SharedReg445_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg445_out;
SharedReg988_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg988_out;
SharedReg1053_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1053_out;
SharedReg746_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg746_out;
SharedReg1116_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1116_out;
   MUX_Product50_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1117_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg42_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg746_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1116_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg986_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg878_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1012_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg577_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg678_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg445_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg988_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1053_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product50_2_impl_1_out);

   Delay1No417_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product50_2_impl_1_out,
                 Y => Delay1No417_out);

Delay1No418_out_to_Product50_3_impl_parent_implementedSystem_port_0_cast <= Delay1No418_out;
Delay1No419_out_to_Product50_3_impl_parent_implementedSystem_port_1_cast <= Delay1No419_out;
   Product50_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product50_3_impl_out,
                 X => Delay1No418_out_to_Product50_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No419_out_to_Product50_3_impl_parent_implementedSystem_port_1_cast);

SharedReg176_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg176_out;
SharedReg111_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg111_out;
SharedReg1106_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1106_out;
SharedReg1148_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1148_out;
SharedReg1113_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1113_out;
SharedReg1129_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1129_out;
SharedReg1149_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1149_out;
SharedReg1136_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1136_out;
SharedReg1137_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1137_out;
SharedReg1135_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1135_out;
SharedReg1114_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1114_out;
SharedReg1115_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1115_out;
   MUX_Product50_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg176_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg111_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1114_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1115_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1106_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1148_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1113_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1129_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1149_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1136_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1137_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1135_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product50_3_impl_0_out);

   Delay1No418_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product50_3_impl_0_out,
                 Y => Delay1No418_out);

SharedReg1116_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1116_out;
SharedReg1117_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1117_out;
SharedReg199_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg199_out;
SharedReg990_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg990_out;
SharedReg792_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg792_out;
SharedReg1017_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1017_out;
SharedReg581_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg581_out;
SharedReg683_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg683_out;
SharedReg580_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg580_out;
SharedReg1020_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1020_out;
SharedReg1059_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1059_out;
SharedReg451_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg451_out;
   MUX_Product50_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1116_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1117_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1059_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg451_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg199_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg990_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg792_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1017_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg581_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg683_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg580_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1020_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product50_3_impl_1_out);

   Delay1No419_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product50_3_impl_1_out,
                 Y => Delay1No419_out);

Delay1No420_out_to_Product50_4_impl_parent_implementedSystem_port_0_cast <= Delay1No420_out;
Delay1No421_out_to_Product50_4_impl_parent_implementedSystem_port_1_cast <= Delay1No421_out;
   Product50_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product50_4_impl_out,
                 X => Delay1No420_out_to_Product50_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No421_out_to_Product50_4_impl_parent_implementedSystem_port_1_cast);

SharedReg1114_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1114_out;
SharedReg1115_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1115_out;
SharedReg53_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg53_out;
SharedReg115_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg115_out;
SharedReg1106_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1106_out;
SharedReg1148_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1148_out;
SharedReg1113_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1113_out;
SharedReg1129_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1129_out;
SharedReg1149_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1149_out;
SharedReg1136_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1136_out;
SharedReg1137_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1137_out;
SharedReg1135_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1135_out;
   MUX_Product50_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1114_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1115_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1137_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1135_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg53_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg115_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1106_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1148_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1113_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1129_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1149_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1136_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product50_4_impl_0_out);

   Delay1No420_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product50_4_impl_0_out,
                 Y => Delay1No420_out);

SharedReg1026_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1026_out;
SharedReg705_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg705_out;
SharedReg1116_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1116_out;
SharedReg1117_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1117_out;
SharedReg177_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg177_out;
SharedReg865_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg865_out;
SharedReg797_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg797_out;
SharedReg1022_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1022_out;
SharedReg585_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg585_out;
SharedReg689_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg689_out;
SharedReg458_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg458_out;
SharedReg1024_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1024_out;
   MUX_Product50_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1026_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg705_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg458_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1024_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1116_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1117_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg177_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg865_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg797_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1022_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg585_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg689_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product50_4_impl_1_out);

   Delay1No421_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product50_4_impl_1_out,
                 Y => Delay1No421_out);

Delay1No422_out_to_Product50_5_impl_parent_implementedSystem_port_0_cast <= Delay1No422_out;
Delay1No423_out_to_Product50_5_impl_parent_implementedSystem_port_1_cast <= Delay1No423_out;
   Product50_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product50_5_impl_out,
                 X => Delay1No422_out_to_Product50_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No423_out_to_Product50_5_impl_parent_implementedSystem_port_1_cast);

SharedReg1137_out_to_MUX_Product50_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1137_out;
SharedReg1135_out_to_MUX_Product50_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1135_out;
SharedReg1114_out_to_MUX_Product50_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1114_out;
SharedReg1115_out_to_MUX_Product50_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1115_out;
SharedReg314_out_to_MUX_Product50_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg314_out;
SharedReg151_out_to_MUX_Product50_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg151_out;
SharedReg1106_out_to_MUX_Product50_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1106_out;
SharedReg1148_out_to_MUX_Product50_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1148_out;
SharedReg1113_out_to_MUX_Product50_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1113_out;
SharedReg1129_out_to_MUX_Product50_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1129_out;
SharedReg1149_out_to_MUX_Product50_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1149_out;
SharedReg1136_out_to_MUX_Product50_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1136_out;
   MUX_Product50_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1137_out_to_MUX_Product50_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1135_out_to_MUX_Product50_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1149_out_to_MUX_Product50_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1136_out_to_MUX_Product50_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1114_out_to_MUX_Product50_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1115_out_to_MUX_Product50_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg314_out_to_MUX_Product50_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg151_out_to_MUX_Product50_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1106_out_to_MUX_Product50_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1148_out_to_MUX_Product50_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1113_out_to_MUX_Product50_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1129_out_to_MUX_Product50_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product50_5_impl_0_out);

   Delay1No422_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product50_5_impl_0_out,
                 Y => Delay1No422_out);

SharedReg464_out_to_MUX_Product50_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg464_out;
SharedReg1031_out_to_MUX_Product50_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1031_out;
SharedReg1064_out_to_MUX_Product50_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1064_out;
SharedReg764_out_to_MUX_Product50_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg764_out;
SharedReg1116_out_to_MUX_Product50_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1116_out;
SharedReg1117_out_to_MUX_Product50_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1117_out;
SharedReg54_out_to_MUX_Product50_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg54_out;
SharedReg997_out_to_MUX_Product50_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg997_out;
SharedReg772_out_to_MUX_Product50_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg772_out;
SharedReg1060_out_to_MUX_Product50_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1060_out;
SharedReg695_out_to_MUX_Product50_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg695_out;
SharedReg868_out_to_MUX_Product50_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg868_out;
   MUX_Product50_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg464_out_to_MUX_Product50_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1031_out_to_MUX_Product50_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg695_out_to_MUX_Product50_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg868_out_to_MUX_Product50_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1064_out_to_MUX_Product50_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg764_out_to_MUX_Product50_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1116_out_to_MUX_Product50_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1117_out_to_MUX_Product50_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg54_out_to_MUX_Product50_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg997_out_to_MUX_Product50_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg772_out_to_MUX_Product50_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1060_out_to_MUX_Product50_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product50_5_impl_1_out);

   Delay1No423_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product50_5_impl_1_out,
                 Y => Delay1No423_out);

Delay1No424_out_to_Product50_6_impl_parent_implementedSystem_port_0_cast <= Delay1No424_out;
Delay1No425_out_to_Product50_6_impl_parent_implementedSystem_port_1_cast <= Delay1No425_out;
   Product50_6_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product50_6_impl_out,
                 X => Delay1No424_out_to_Product50_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No425_out_to_Product50_6_impl_parent_implementedSystem_port_1_cast);

SharedReg1136_out_to_MUX_Product50_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1136_out;
SharedReg1137_out_to_MUX_Product50_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1137_out;
SharedReg1135_out_to_MUX_Product50_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1135_out;
SharedReg1114_out_to_MUX_Product50_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1114_out;
SharedReg1115_out_to_MUX_Product50_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1115_out;
SharedReg382_out_to_MUX_Product50_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg382_out;
SharedReg124_out_to_MUX_Product50_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg124_out;
SharedReg1106_out_to_MUX_Product50_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1106_out;
SharedReg1148_out_to_MUX_Product50_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1148_out;
SharedReg1113_out_to_MUX_Product50_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1113_out;
SharedReg1129_out_to_MUX_Product50_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1129_out;
SharedReg1149_out_to_MUX_Product50_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1149_out;
   MUX_Product50_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1136_out_to_MUX_Product50_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1137_out_to_MUX_Product50_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1129_out_to_MUX_Product50_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1149_out_to_MUX_Product50_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1135_out_to_MUX_Product50_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1114_out_to_MUX_Product50_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1115_out_to_MUX_Product50_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg382_out_to_MUX_Product50_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg124_out_to_MUX_Product50_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1106_out_to_MUX_Product50_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1148_out_to_MUX_Product50_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1113_out_to_MUX_Product50_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product50_6_impl_0_out);

   Delay1No424_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product50_6_impl_0_out,
                 Y => Delay1No424_out);

SharedReg871_out_to_MUX_Product50_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg871_out;
SharedReg699_out_to_MUX_Product50_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg699_out;
SharedReg1078_out_to_MUX_Product50_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1078_out;
SharedReg1079_out_to_MUX_Product50_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1079_out;
SharedReg473_out_to_MUX_Product50_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg473_out;
SharedReg1116_out_to_MUX_Product50_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1116_out;
SharedReg1117_out_to_MUX_Product50_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1117_out;
SharedReg226_out_to_MUX_Product50_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg226_out;
SharedReg1066_out_to_MUX_Product50_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1066_out;
SharedReg1090_out_to_MUX_Product50_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1090_out;
SharedReg1075_out_to_MUX_Product50_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1075_out;
SharedReg872_out_to_MUX_Product50_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg872_out;
   MUX_Product50_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg871_out_to_MUX_Product50_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg699_out_to_MUX_Product50_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1075_out_to_MUX_Product50_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg872_out_to_MUX_Product50_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1078_out_to_MUX_Product50_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1079_out_to_MUX_Product50_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg473_out_to_MUX_Product50_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1116_out_to_MUX_Product50_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1117_out_to_MUX_Product50_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg226_out_to_MUX_Product50_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1066_out_to_MUX_Product50_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1090_out_to_MUX_Product50_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product50_6_impl_1_out);

   Delay1No425_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product50_6_impl_1_out,
                 Y => Delay1No425_out);

Delay1No426_out_to_Product122_0_impl_parent_implementedSystem_port_0_cast <= Delay1No426_out;
Delay1No427_out_to_Product122_0_impl_parent_implementedSystem_port_1_cast <= Delay1No427_out;
   Product122_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product122_0_impl_out,
                 X => Delay1No426_out_to_Product122_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No427_out_to_Product122_0_impl_parent_implementedSystem_port_1_cast);

SharedReg1129_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1129_out;
SharedReg1149_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1149_out;
SharedReg1136_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1136_out;
SharedReg1137_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1137_out;
SharedReg1135_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1135_out;
SharedReg1114_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1114_out;
SharedReg564_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg564_out;
SharedReg1104_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1104_out;
SharedReg1117_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1117_out;
SharedReg1118_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1118_out;
SharedReg1148_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1148_out;
SharedReg1113_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1113_out;
   MUX_Product122_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1129_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1149_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1148_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1113_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1136_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1137_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1135_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1114_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg564_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1104_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1117_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1118_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product122_0_impl_0_out);

   Delay1No426_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product122_0_impl_0_out,
                 Y => Delay1No426_out);

SharedReg1094_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1094_out;
SharedReg1004_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1004_out;
SharedReg981_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg981_out;
SharedReg666_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg666_out;
SharedReg1073_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1073_out;
SharedReg1095_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1095_out;
SharedReg1115_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1115_out;
SharedReg565_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg565_out;
SharedReg250_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg250_out;
SharedReg34_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg34_out;
SharedReg1070_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1070_out;
SharedReg778_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg778_out;
   MUX_Product122_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1094_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1004_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1070_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg778_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg981_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg666_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1073_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1095_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1115_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg565_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg250_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg34_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product122_0_impl_1_out);

   Delay1No427_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product122_0_impl_1_out,
                 Y => Delay1No427_out);

Delay1No428_out_to_Product122_1_impl_parent_implementedSystem_port_0_cast <= Delay1No428_out;
Delay1No429_out_to_Product122_1_impl_parent_implementedSystem_port_1_cast <= Delay1No429_out;
   Product122_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product122_1_impl_out,
                 X => Delay1No428_out_to_Product122_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No429_out_to_Product122_1_impl_parent_implementedSystem_port_1_cast);

SharedReg1148_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1148_out;
SharedReg1113_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1113_out;
SharedReg1129_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1129_out;
SharedReg1149_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1149_out;
SharedReg1136_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1136_out;
SharedReg1137_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1137_out;
SharedReg1135_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1135_out;
SharedReg1114_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1114_out;
SharedReg570_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg570_out;
SharedReg1104_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1104_out;
SharedReg1117_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1117_out;
SharedReg1118_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1118_out;
   MUX_Product122_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1148_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1113_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1117_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1118_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1129_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1149_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1136_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1137_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1135_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1114_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg570_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1104_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product122_1_impl_0_out);

   Delay1No428_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product122_1_impl_0_out,
                 Y => Delay1No428_out);

SharedReg1042_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1042_out;
SharedReg786_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg786_out;
SharedReg1081_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1081_out;
SharedReg984_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg984_out;
SharedReg854_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg854_out;
SharedReg570_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg570_out;
SharedReg1045_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1045_out;
SharedReg784_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg784_out;
SharedReg1115_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1115_out;
SharedReg571_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg571_out;
SharedReg255_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg255_out;
SharedReg39_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg39_out;
   MUX_Product122_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1042_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg786_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg255_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg39_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1081_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg984_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg854_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg570_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1045_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg784_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1115_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg571_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product122_1_impl_1_out);

   Delay1No429_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product122_1_impl_1_out,
                 Y => Delay1No429_out);

Delay1No430_out_to_Product122_2_impl_parent_implementedSystem_port_0_cast <= Delay1No430_out;
Delay1No431_out_to_Product122_2_impl_parent_implementedSystem_port_1_cast <= Delay1No431_out;
   Product122_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product122_2_impl_out,
                 X => Delay1No430_out_to_Product122_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No431_out_to_Product122_2_impl_parent_implementedSystem_port_1_cast);

SharedReg1117_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1117_out;
SharedReg1118_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1118_out;
SharedReg1148_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1148_out;
SharedReg1113_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1113_out;
SharedReg1129_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1129_out;
SharedReg1149_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1149_out;
SharedReg1136_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1136_out;
SharedReg1137_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1137_out;
SharedReg1135_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1135_out;
SharedReg1114_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1114_out;
SharedReg445_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg445_out;
SharedReg1104_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1104_out;
   MUX_Product122_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1117_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1118_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg445_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1104_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1148_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1113_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1129_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1149_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1136_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1137_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1135_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1114_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product122_2_impl_0_out);

   Delay1No430_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product122_2_impl_0_out,
                 Y => Delay1No430_out);

SharedReg261_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg261_out;
SharedReg42_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg42_out;
SharedReg1012_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1012_out;
SharedReg879_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg879_out;
SharedReg1047_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1047_out;
SharedReg858_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg858_out;
SharedReg858_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg858_out;
SharedReg576_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg576_out;
SharedReg1015_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1015_out;
SharedReg754_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg754_out;
SharedReg1115_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1115_out;
SharedReg446_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg446_out;
   MUX_Product122_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg261_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg42_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1115_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg446_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1012_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg879_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1047_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg858_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg858_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg576_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1015_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg754_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product122_2_impl_1_out);

   Delay1No431_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product122_2_impl_1_out,
                 Y => Delay1No431_out);

Delay1No432_out_to_Product122_3_impl_parent_implementedSystem_port_0_cast <= Delay1No432_out;
Delay1No433_out_to_Product122_3_impl_parent_implementedSystem_port_1_cast <= Delay1No433_out;
   Product122_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product122_3_impl_out,
                 X => Delay1No432_out_to_Product122_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No433_out_to_Product122_3_impl_parent_implementedSystem_port_1_cast);

SharedReg1104_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1104_out;
SharedReg1117_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1117_out;
SharedReg1118_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1118_out;
SharedReg1148_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1148_out;
SharedReg1113_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1113_out;
SharedReg1129_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1129_out;
SharedReg1149_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1149_out;
SharedReg1136_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1136_out;
SharedReg1137_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1137_out;
SharedReg1135_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1135_out;
SharedReg1114_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1114_out;
SharedReg580_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg580_out;
   MUX_Product122_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1104_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1117_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1114_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg580_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1118_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1148_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1113_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1129_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1149_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1136_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1137_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1135_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product122_3_impl_0_out);

   Delay1No432_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product122_3_impl_0_out,
                 Y => Delay1No432_out);

SharedReg581_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg581_out;
SharedReg245_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg245_out;
SharedReg199_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg199_out;
SharedReg1017_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1017_out;
SharedReg760_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg760_out;
SharedReg1054_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1054_out;
SharedReg990_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg990_out;
SharedReg861_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg861_out;
SharedReg683_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg683_out;
SharedReg1056_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1056_out;
SharedReg759_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg759_out;
SharedReg1115_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1115_out;
   MUX_Product122_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg581_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg245_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg759_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1115_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg199_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1017_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg760_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1054_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg990_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg861_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg683_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1056_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product122_3_impl_1_out);

   Delay1No433_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product122_3_impl_1_out,
                 Y => Delay1No433_out);

Delay1No434_out_to_Product122_4_impl_parent_implementedSystem_port_0_cast <= Delay1No434_out;
Delay1No435_out_to_Product122_4_impl_parent_implementedSystem_port_1_cast <= Delay1No435_out;
   Product122_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product122_4_impl_out,
                 X => Delay1No434_out_to_Product122_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No435_out_to_Product122_4_impl_parent_implementedSystem_port_1_cast);

SharedReg1114_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1114_out;
SharedReg458_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg458_out;
SharedReg1104_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1104_out;
SharedReg1117_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1117_out;
SharedReg1118_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1118_out;
SharedReg1148_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1148_out;
SharedReg1113_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1113_out;
SharedReg1129_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1129_out;
SharedReg1149_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1149_out;
SharedReg1136_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1136_out;
SharedReg1137_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1137_out;
SharedReg1135_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1135_out;
   MUX_Product122_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1114_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg458_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1137_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1135_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1104_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1117_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1118_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1148_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1113_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1129_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1149_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1136_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product122_4_impl_0_out);

   Delay1No434_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product122_4_impl_0_out,
                 Y => Delay1No434_out);

SharedReg713_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg713_out;
SharedReg1115_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1115_out;
SharedReg459_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg459_out;
SharedReg207_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg207_out;
SharedReg177_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg177_out;
SharedReg993_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg993_out;
SharedReg798_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg798_out;
SharedReg795_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg795_out;
SharedReg993_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg993_out;
SharedReg865_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg865_out;
SharedReg584_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg584_out;
SharedReg798_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg798_out;
   MUX_Product122_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg713_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1115_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg584_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg798_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg459_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg207_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg177_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg993_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg798_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg795_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg993_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg865_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product122_4_impl_1_out);

   Delay1No435_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product122_4_impl_1_out,
                 Y => Delay1No435_out);

Delay1No436_out_to_Product122_5_impl_parent_implementedSystem_port_0_cast <= Delay1No436_out;
Delay1No437_out_to_Product122_5_impl_parent_implementedSystem_port_1_cast <= Delay1No437_out;
   Product122_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product122_5_impl_out,
                 X => Delay1No436_out_to_Product122_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No437_out_to_Product122_5_impl_parent_implementedSystem_port_1_cast);

SharedReg1137_out_to_MUX_Product122_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1137_out;
SharedReg1135_out_to_MUX_Product122_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1135_out;
SharedReg1114_out_to_MUX_Product122_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1114_out;
SharedReg712_out_to_MUX_Product122_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg712_out;
SharedReg1104_out_to_MUX_Product122_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1104_out;
SharedReg1117_out_to_MUX_Product122_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1117_out;
SharedReg1118_out_to_MUX_Product122_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1118_out;
SharedReg1148_out_to_MUX_Product122_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1148_out;
SharedReg1113_out_to_MUX_Product122_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1113_out;
SharedReg1129_out_to_MUX_Product122_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1129_out;
SharedReg1149_out_to_MUX_Product122_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1149_out;
SharedReg1136_out_to_MUX_Product122_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1136_out;
   MUX_Product122_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1137_out_to_MUX_Product122_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1135_out_to_MUX_Product122_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1149_out_to_MUX_Product122_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1136_out_to_MUX_Product122_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1114_out_to_MUX_Product122_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg712_out_to_MUX_Product122_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1104_out_to_MUX_Product122_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1117_out_to_MUX_Product122_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1118_out_to_MUX_Product122_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1148_out_to_MUX_Product122_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1113_out_to_MUX_Product122_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1129_out_to_MUX_Product122_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product122_5_impl_0_out);

   Delay1No436_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product122_5_impl_0_out,
                 Y => Delay1No436_out);

SharedReg589_out_to_MUX_Product122_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg589_out;
SharedReg1062_out_to_MUX_Product122_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1062_out;
SharedReg474_out_to_MUX_Product122_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg474_out;
SharedReg1115_out_to_MUX_Product122_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1115_out;
SharedReg713_out_to_MUX_Product122_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg713_out;
SharedReg213_out_to_MUX_Product122_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg213_out;
SharedReg54_out_to_MUX_Product122_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg54_out;
SharedReg1028_out_to_MUX_Product122_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1028_out;
SharedReg1062_out_to_MUX_Product122_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1062_out;
SharedReg770_out_to_MUX_Product122_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg770_out;
SharedReg997_out_to_MUX_Product122_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg997_out;
SharedReg997_out_to_MUX_Product122_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg997_out;
   MUX_Product122_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg589_out_to_MUX_Product122_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1062_out_to_MUX_Product122_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg997_out_to_MUX_Product122_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg997_out_to_MUX_Product122_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg474_out_to_MUX_Product122_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1115_out_to_MUX_Product122_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg713_out_to_MUX_Product122_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg213_out_to_MUX_Product122_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg54_out_to_MUX_Product122_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1028_out_to_MUX_Product122_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1062_out_to_MUX_Product122_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg770_out_to_MUX_Product122_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product122_5_impl_1_out);

   Delay1No437_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product122_5_impl_1_out,
                 Y => Delay1No437_out);

Delay1No438_out_to_Product122_6_impl_parent_implementedSystem_port_0_cast <= Delay1No438_out;
Delay1No439_out_to_Product122_6_impl_parent_implementedSystem_port_1_cast <= Delay1No439_out;
   Product122_6_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product122_6_impl_out,
                 X => Delay1No438_out_to_Product122_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No439_out_to_Product122_6_impl_parent_implementedSystem_port_1_cast);

SharedReg1136_out_to_MUX_Product122_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1136_out;
SharedReg1137_out_to_MUX_Product122_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1137_out;
SharedReg1135_out_to_MUX_Product122_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1135_out;
SharedReg1114_out_to_MUX_Product122_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1114_out;
SharedReg595_out_to_MUX_Product122_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg595_out;
SharedReg1104_out_to_MUX_Product122_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1104_out;
SharedReg1117_out_to_MUX_Product122_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1117_out;
SharedReg1118_out_to_MUX_Product122_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1118_out;
SharedReg1148_out_to_MUX_Product122_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1148_out;
SharedReg1113_out_to_MUX_Product122_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1113_out;
SharedReg1129_out_to_MUX_Product122_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1129_out;
SharedReg1149_out_to_MUX_Product122_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1149_out;
   MUX_Product122_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1136_out_to_MUX_Product122_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1137_out_to_MUX_Product122_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1129_out_to_MUX_Product122_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1149_out_to_MUX_Product122_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1135_out_to_MUX_Product122_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1114_out_to_MUX_Product122_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg595_out_to_MUX_Product122_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1104_out_to_MUX_Product122_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1117_out_to_MUX_Product122_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1118_out_to_MUX_Product122_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1148_out_to_MUX_Product122_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1113_out_to_MUX_Product122_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product122_6_impl_0_out);

   Delay1No438_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product122_6_impl_0_out,
                 Y => Delay1No438_out);

SharedReg1001_out_to_MUX_Product122_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1001_out;
SharedReg871_out_to_MUX_Product122_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg871_out;
SharedReg1091_out_to_MUX_Product122_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1091_out;
SharedReg1089_out_to_MUX_Product122_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1089_out;
SharedReg1115_out_to_MUX_Product122_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1115_out;
SharedReg596_out_to_MUX_Product122_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg596_out;
SharedReg188_out_to_MUX_Product122_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg188_out;
SharedReg226_out_to_MUX_Product122_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg226_out;
SharedReg1075_out_to_MUX_Product122_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1075_out;
SharedReg1102_out_to_MUX_Product122_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1102_out;
SharedReg1088_out_to_MUX_Product122_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1088_out;
SharedReg1066_out_to_MUX_Product122_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1066_out;
   MUX_Product122_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1001_out_to_MUX_Product122_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg871_out_to_MUX_Product122_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1088_out_to_MUX_Product122_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1066_out_to_MUX_Product122_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1091_out_to_MUX_Product122_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1089_out_to_MUX_Product122_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1115_out_to_MUX_Product122_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg596_out_to_MUX_Product122_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg188_out_to_MUX_Product122_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg226_out_to_MUX_Product122_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1075_out_to_MUX_Product122_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1102_out_to_MUX_Product122_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product122_6_impl_1_out);

   Delay1No439_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product122_6_impl_1_out,
                 Y => Delay1No439_out);

Delay1No440_out_to_Product221_0_impl_parent_implementedSystem_port_0_cast <= Delay1No440_out;
Delay1No441_out_to_Product221_0_impl_parent_implementedSystem_port_1_cast <= Delay1No441_out;
   Product221_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product221_0_impl_out,
                 X => Delay1No440_out_to_Product221_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No441_out_to_Product221_0_impl_parent_implementedSystem_port_1_cast);

SharedReg1131_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1131_out;
SharedReg1153_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1153_out;
SharedReg1140_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1140_out;
SharedReg1141_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1141_out;
SharedReg1139_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1139_out;
SharedReg1126_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1126_out;
SharedReg1158_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1158_out;
SharedReg1159_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1159_out;
SharedReg160_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg160_out;
SharedReg1106_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1106_out;
SharedReg1152_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1152_out;
SharedReg1125_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1125_out;
   MUX_Product221_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1131_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1153_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1152_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1125_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1140_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1141_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1139_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1126_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1158_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1159_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg160_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1106_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product221_0_impl_0_out);

   Delay1No440_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product221_0_impl_0_out,
                 Y => Delay1No440_out);

SharedReg1070_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1070_out;
SharedReg850_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg850_out;
SharedReg849_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg849_out;
SharedReg564_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg564_out;
SharedReg1040_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1040_out;
SharedReg1100_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1100_out;
SharedReg666_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg666_out;
SharedReg667_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg667_out;
SharedReg1117_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1117_out;
SharedReg251_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg251_out;
SharedReg1037_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1037_out;
SharedReg777_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg777_out;
   MUX_Product221_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1070_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg850_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1037_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg777_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg849_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg564_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1040_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1100_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg666_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg667_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1117_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg251_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product221_0_impl_1_out);

   Delay1No441_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product221_0_impl_1_out,
                 Y => Delay1No441_out);

Delay1No442_out_to_Product221_1_impl_parent_implementedSystem_port_0_cast <= Delay1No442_out;
Delay1No443_out_to_Product221_1_impl_parent_implementedSystem_port_1_cast <= Delay1No443_out;
   Product221_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product221_1_impl_out,
                 X => Delay1No442_out_to_Product221_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No443_out_to_Product221_1_impl_parent_implementedSystem_port_1_cast);

SharedReg1152_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1152_out;
SharedReg1125_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1125_out;
SharedReg1131_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1131_out;
SharedReg1153_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1153_out;
SharedReg1140_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1140_out;
SharedReg1141_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1141_out;
SharedReg1139_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1139_out;
SharedReg1126_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1126_out;
SharedReg1158_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1158_out;
SharedReg1159_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1159_out;
SharedReg42_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg42_out;
SharedReg1106_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1106_out;
   MUX_Product221_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1152_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1125_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg42_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1106_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1131_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1153_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1140_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1141_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1139_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1126_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1158_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1159_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product221_1_impl_0_out);

   Delay1No442_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product221_1_impl_0_out,
                 Y => Delay1No442_out);

SharedReg1007_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1007_out;
SharedReg785_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg785_out;
SharedReg1042_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1042_out;
SharedReg673_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg673_out;
SharedReg672_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg672_out;
SharedReg438_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg438_out;
SharedReg1010_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1010_out;
SharedReg1087_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1087_out;
SharedReg672_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg672_out;
SharedReg673_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg673_out;
SharedReg1117_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1117_out;
SharedReg256_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg256_out;
   MUX_Product221_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1007_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg785_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1117_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg256_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1042_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg673_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg672_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg438_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1010_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1087_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg672_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg673_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product221_1_impl_1_out);

   Delay1No443_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product221_1_impl_1_out,
                 Y => Delay1No443_out);

Delay1No444_out_to_Product221_2_impl_parent_implementedSystem_port_0_cast <= Delay1No444_out;
Delay1No445_out_to_Product221_2_impl_parent_implementedSystem_port_1_cast <= Delay1No445_out;
   Product221_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product221_2_impl_out,
                 X => Delay1No444_out_to_Product221_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No445_out_to_Product221_2_impl_parent_implementedSystem_port_1_cast);

SharedReg199_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg199_out;
SharedReg1106_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1106_out;
SharedReg1152_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1152_out;
SharedReg1125_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1125_out;
SharedReg1131_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1131_out;
SharedReg1153_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1153_out;
SharedReg1140_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1140_out;
SharedReg1141_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1141_out;
SharedReg1139_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1139_out;
SharedReg1126_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1126_out;
SharedReg1158_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1158_out;
SharedReg1159_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1159_out;
   MUX_Product221_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg199_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1106_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1158_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1159_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1152_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1125_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1131_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1153_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1140_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1141_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1139_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1126_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product221_2_impl_0_out);

   Delay1No444_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product221_2_impl_0_out,
                 Y => Delay1No444_out);

SharedReg1117_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1117_out;
SharedReg262_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg262_out;
SharedReg986_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg986_out;
SharedReg878_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg878_out;
SharedReg1012_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1012_out;
SharedReg577_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg577_out;
SharedReg678_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg678_out;
SharedReg445_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg445_out;
SharedReg988_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg988_out;
SharedReg1053_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1053_out;
SharedReg576_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg576_out;
SharedReg577_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg577_out;
   MUX_Product221_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1117_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg262_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg576_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg577_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg986_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg878_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1012_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg577_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg678_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg445_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg988_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1053_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product221_2_impl_1_out);

   Delay1No445_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product221_2_impl_1_out,
                 Y => Delay1No445_out);

Delay1No446_out_to_Product221_3_impl_parent_implementedSystem_port_0_cast <= Delay1No446_out;
Delay1No447_out_to_Product221_3_impl_parent_implementedSystem_port_1_cast <= Delay1No447_out;
   Product221_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product221_3_impl_out,
                 X => Delay1No446_out_to_Product221_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No447_out_to_Product221_3_impl_parent_implementedSystem_port_1_cast);

SharedReg1159_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1159_out;
SharedReg50_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg50_out;
SharedReg1106_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1106_out;
SharedReg1152_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1152_out;
SharedReg1125_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1125_out;
SharedReg1131_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1131_out;
SharedReg1153_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1153_out;
SharedReg1140_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1140_out;
SharedReg1141_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1141_out;
SharedReg1139_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1139_out;
SharedReg1126_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1126_out;
SharedReg1158_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1158_out;
   MUX_Product221_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1159_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg50_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1126_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1158_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1106_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1152_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1125_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1131_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1153_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1140_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1141_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1139_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product221_3_impl_0_out);

   Delay1No446_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product221_3_impl_0_out,
                 Y => Delay1No446_out);

SharedReg684_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg684_out;
SharedReg1117_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1117_out;
SharedReg246_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg246_out;
SharedReg990_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg990_out;
SharedReg792_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg792_out;
SharedReg1017_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1017_out;
SharedReg581_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg581_out;
SharedReg683_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg683_out;
SharedReg580_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg580_out;
SharedReg1020_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1020_out;
SharedReg1059_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1059_out;
SharedReg683_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg683_out;
   MUX_Product221_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg684_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1117_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1059_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg683_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg246_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg990_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg792_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1017_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg581_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg683_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg580_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1020_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product221_3_impl_1_out);

   Delay1No447_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product221_3_impl_1_out,
                 Y => Delay1No447_out);

Delay1No448_out_to_Product221_4_impl_parent_implementedSystem_port_0_cast <= Delay1No448_out;
Delay1No449_out_to_Product221_4_impl_parent_implementedSystem_port_1_cast <= Delay1No449_out;
   Product221_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product221_4_impl_out,
                 X => Delay1No448_out_to_Product221_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No449_out_to_Product221_4_impl_parent_implementedSystem_port_1_cast);

SharedReg1126_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1126_out;
SharedReg1158_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1158_out;
SharedReg1159_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1159_out;
SharedReg88_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg88_out;
SharedReg1106_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1106_out;
SharedReg1152_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1152_out;
SharedReg1125_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1125_out;
SharedReg1131_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1131_out;
SharedReg1153_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1153_out;
SharedReg1140_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1140_out;
SharedReg1141_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1141_out;
SharedReg1139_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1139_out;
   MUX_Product221_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1126_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1158_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1141_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1139_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1159_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg88_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1106_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1152_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1125_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1131_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1153_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1140_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product221_4_impl_0_out);

   Delay1No448_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product221_4_impl_0_out,
                 Y => Delay1No448_out);

SharedReg1026_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1026_out;
SharedReg584_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg584_out;
SharedReg585_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg585_out;
SharedReg1117_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1117_out;
SharedReg208_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg208_out;
SharedReg865_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg865_out;
SharedReg797_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg797_out;
SharedReg1022_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1022_out;
SharedReg585_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg585_out;
SharedReg689_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg689_out;
SharedReg458_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg458_out;
SharedReg1024_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1024_out;
   MUX_Product221_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1026_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg584_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg458_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1024_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg585_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1117_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg208_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg865_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg797_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1022_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg585_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg689_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product221_4_impl_1_out);

   Delay1No449_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product221_4_impl_1_out,
                 Y => Delay1No449_out);

Delay1No450_out_to_Product221_5_impl_parent_implementedSystem_port_0_cast <= Delay1No450_out;
Delay1No451_out_to_Product221_5_impl_parent_implementedSystem_port_1_cast <= Delay1No451_out;
   Product221_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product221_5_impl_out,
                 X => Delay1No450_out_to_Product221_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No451_out_to_Product221_5_impl_parent_implementedSystem_port_1_cast);

SharedReg1141_out_to_MUX_Product221_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1141_out;
SharedReg1139_out_to_MUX_Product221_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1139_out;
SharedReg1126_out_to_MUX_Product221_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1126_out;
SharedReg1158_out_to_MUX_Product221_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1158_out;
SharedReg1159_out_to_MUX_Product221_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1159_out;
SharedReg226_out_to_MUX_Product221_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg226_out;
SharedReg1106_out_to_MUX_Product221_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1106_out;
SharedReg1152_out_to_MUX_Product221_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1152_out;
SharedReg1125_out_to_MUX_Product221_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1125_out;
SharedReg1131_out_to_MUX_Product221_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1131_out;
SharedReg1153_out_to_MUX_Product221_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1153_out;
SharedReg1140_out_to_MUX_Product221_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1140_out;
   MUX_Product221_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1141_out_to_MUX_Product221_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1139_out_to_MUX_Product221_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1153_out_to_MUX_Product221_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1140_out_to_MUX_Product221_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1126_out_to_MUX_Product221_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1158_out_to_MUX_Product221_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1159_out_to_MUX_Product221_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg226_out_to_MUX_Product221_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1106_out_to_MUX_Product221_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1152_out_to_MUX_Product221_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1125_out_to_MUX_Product221_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1131_out_to_MUX_Product221_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product221_5_impl_0_out);

   Delay1No450_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product221_5_impl_0_out,
                 Y => Delay1No450_out);

SharedReg464_out_to_MUX_Product221_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg464_out;
SharedReg1031_out_to_MUX_Product221_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1031_out;
SharedReg1064_out_to_MUX_Product221_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1064_out;
SharedReg464_out_to_MUX_Product221_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg464_out;
SharedReg465_out_to_MUX_Product221_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg465_out;
SharedReg1117_out_to_MUX_Product221_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1117_out;
SharedReg214_out_to_MUX_Product221_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg214_out;
SharedReg997_out_to_MUX_Product221_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg997_out;
SharedReg772_out_to_MUX_Product221_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg772_out;
SharedReg1060_out_to_MUX_Product221_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1060_out;
SharedReg695_out_to_MUX_Product221_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg695_out;
SharedReg868_out_to_MUX_Product221_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg868_out;
   MUX_Product221_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg464_out_to_MUX_Product221_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1031_out_to_MUX_Product221_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg695_out_to_MUX_Product221_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg868_out_to_MUX_Product221_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1064_out_to_MUX_Product221_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg464_out_to_MUX_Product221_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg465_out_to_MUX_Product221_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1117_out_to_MUX_Product221_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg214_out_to_MUX_Product221_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg997_out_to_MUX_Product221_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg772_out_to_MUX_Product221_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1060_out_to_MUX_Product221_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product221_5_impl_1_out);

   Delay1No451_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product221_5_impl_1_out,
                 Y => Delay1No451_out);

Delay1No452_out_to_Product221_6_impl_parent_implementedSystem_port_0_cast <= Delay1No452_out;
Delay1No453_out_to_Product221_6_impl_parent_implementedSystem_port_1_cast <= Delay1No453_out;
   Product221_6_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product221_6_impl_out,
                 X => Delay1No452_out_to_Product221_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No453_out_to_Product221_6_impl_parent_implementedSystem_port_1_cast);

SharedReg1140_out_to_MUX_Product221_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1140_out;
SharedReg1141_out_to_MUX_Product221_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1141_out;
SharedReg1139_out_to_MUX_Product221_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1139_out;
SharedReg1126_out_to_MUX_Product221_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1126_out;
SharedReg1158_out_to_MUX_Product221_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1158_out;
SharedReg1159_out_to_MUX_Product221_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1159_out;
SharedReg390_out_to_MUX_Product221_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg390_out;
SharedReg1106_out_to_MUX_Product221_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1106_out;
SharedReg1152_out_to_MUX_Product221_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1152_out;
SharedReg1125_out_to_MUX_Product221_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1125_out;
SharedReg1131_out_to_MUX_Product221_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1131_out;
SharedReg1153_out_to_MUX_Product221_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1153_out;
   MUX_Product221_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1140_out_to_MUX_Product221_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1141_out_to_MUX_Product221_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1131_out_to_MUX_Product221_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1153_out_to_MUX_Product221_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1139_out_to_MUX_Product221_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1126_out_to_MUX_Product221_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1158_out_to_MUX_Product221_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1159_out_to_MUX_Product221_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg390_out_to_MUX_Product221_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1106_out_to_MUX_Product221_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1152_out_to_MUX_Product221_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1125_out_to_MUX_Product221_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product221_6_impl_0_out);

   Delay1No452_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product221_6_impl_0_out,
                 Y => Delay1No452_out);

SharedReg871_out_to_MUX_Product221_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg871_out;
SharedReg699_out_to_MUX_Product221_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg699_out;
SharedReg1078_out_to_MUX_Product221_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1078_out;
SharedReg1079_out_to_MUX_Product221_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1079_out;
SharedReg699_out_to_MUX_Product221_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg699_out;
SharedReg700_out_to_MUX_Product221_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg700_out;
SharedReg1117_out_to_MUX_Product221_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1117_out;
SharedReg189_out_to_MUX_Product221_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg189_out;
SharedReg1066_out_to_MUX_Product221_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1066_out;
SharedReg1090_out_to_MUX_Product221_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1090_out;
SharedReg1075_out_to_MUX_Product221_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1075_out;
SharedReg872_out_to_MUX_Product221_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg872_out;
   MUX_Product221_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg871_out_to_MUX_Product221_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg699_out_to_MUX_Product221_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1075_out_to_MUX_Product221_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg872_out_to_MUX_Product221_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1078_out_to_MUX_Product221_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1079_out_to_MUX_Product221_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg699_out_to_MUX_Product221_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg700_out_to_MUX_Product221_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1117_out_to_MUX_Product221_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg189_out_to_MUX_Product221_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1066_out_to_MUX_Product221_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1090_out_to_MUX_Product221_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product221_6_impl_1_out);

   Delay1No453_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product221_6_impl_1_out,
                 Y => Delay1No453_out);

Delay1No454_out_to_Product321_0_impl_parent_implementedSystem_port_0_cast <= Delay1No454_out;
Delay1No455_out_to_Product321_0_impl_parent_implementedSystem_port_1_cast <= Delay1No455_out;
   Product321_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product321_0_impl_out,
                 X => Delay1No454_out_to_Product321_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No455_out_to_Product321_0_impl_parent_implementedSystem_port_1_cast);

SharedReg1094_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1094_out;
SharedReg1004_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1004_out;
SharedReg981_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg981_out;
SharedReg666_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg666_out;
SharedReg1073_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1073_out;
SharedReg1095_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1095_out;
SharedReg1158_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1158_out;
SharedReg850_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg850_out;
SharedReg1105_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1105_out;
SharedReg1106_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1106_out;
SharedReg1070_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1070_out;
SharedReg778_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg778_out;
   MUX_Product321_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1094_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1004_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1070_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg778_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg981_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg666_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1073_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1095_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1158_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg850_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1105_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1106_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product321_0_impl_0_out);

   Delay1No454_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_0_impl_0_out,
                 Y => Delay1No454_out);

SharedReg1131_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1131_out;
SharedReg1153_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1153_out;
SharedReg1140_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1140_out;
SharedReg1141_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1141_out;
SharedReg1139_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1139_out;
SharedReg1126_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1126_out;
SharedReg849_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg849_out;
SharedReg1159_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1159_out;
SharedReg432_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg432_out;
SharedReg161_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg161_out;
SharedReg1152_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1152_out;
SharedReg1125_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1125_out;
   MUX_Product321_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1131_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1153_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1152_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1125_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1140_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1141_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1139_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1126_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg849_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1159_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg432_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg161_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product321_0_impl_1_out);

   Delay1No455_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_0_impl_1_out,
                 Y => Delay1No455_out);

Delay1No456_out_to_Product321_1_impl_parent_implementedSystem_port_0_cast <= Delay1No456_out;
Delay1No457_out_to_Product321_1_impl_parent_implementedSystem_port_1_cast <= Delay1No457_out;
   Product321_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product321_1_impl_out,
                 X => Delay1No456_out_to_Product321_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No457_out_to_Product321_1_impl_parent_implementedSystem_port_1_cast);

SharedReg1042_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1042_out;
SharedReg786_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg786_out;
SharedReg1081_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1081_out;
SharedReg984_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg984_out;
SharedReg854_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg854_out;
SharedReg570_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg570_out;
SharedReg1045_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1045_out;
SharedReg784_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg784_out;
SharedReg1158_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1158_out;
SharedReg855_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg855_out;
SharedReg1105_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1105_out;
SharedReg1106_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1106_out;
   MUX_Product321_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1042_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg786_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1105_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1106_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1081_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg984_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg854_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg570_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1045_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg784_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1158_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg855_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product321_1_impl_0_out);

   Delay1No456_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_1_impl_0_out,
                 Y => Delay1No456_out);

SharedReg1152_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1152_out;
SharedReg1125_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1125_out;
SharedReg1131_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1131_out;
SharedReg1153_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1153_out;
SharedReg1140_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1140_out;
SharedReg1141_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1141_out;
SharedReg1139_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1139_out;
SharedReg1126_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1126_out;
SharedReg854_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg854_out;
SharedReg1159_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1159_out;
SharedReg439_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg439_out;
SharedReg43_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg43_out;
   MUX_Product321_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1152_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1125_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg439_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg43_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1131_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1153_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1140_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1141_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1139_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1126_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg854_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1159_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product321_1_impl_1_out);

   Delay1No457_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_1_impl_1_out,
                 Y => Delay1No457_out);

Delay1No458_out_to_Product321_2_impl_parent_implementedSystem_port_0_cast <= Delay1No458_out;
Delay1No459_out_to_Product321_2_impl_parent_implementedSystem_port_1_cast <= Delay1No459_out;
   Product321_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product321_2_impl_out,
                 X => Delay1No458_out_to_Product321_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No459_out_to_Product321_2_impl_parent_implementedSystem_port_1_cast);

SharedReg1105_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1105_out;
SharedReg1106_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1106_out;
SharedReg1012_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1012_out;
SharedReg879_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg879_out;
SharedReg1047_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1047_out;
SharedReg858_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg858_out;
SharedReg858_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg858_out;
SharedReg576_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg576_out;
SharedReg1015_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1015_out;
SharedReg754_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg754_out;
SharedReg1158_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1158_out;
SharedReg679_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg679_out;
   MUX_Product321_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1105_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1106_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1158_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg679_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1012_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg879_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1047_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg858_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg858_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg576_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1015_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg754_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product321_2_impl_0_out);

   Delay1No458_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_2_impl_0_out,
                 Y => Delay1No458_out);

SharedReg747_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg747_out;
SharedReg200_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg200_out;
SharedReg1152_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1152_out;
SharedReg1125_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1125_out;
SharedReg1131_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1131_out;
SharedReg1153_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1153_out;
SharedReg1140_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1140_out;
SharedReg1141_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1141_out;
SharedReg1139_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1139_out;
SharedReg1126_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1126_out;
SharedReg678_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg678_out;
SharedReg1159_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1159_out;
   MUX_Product321_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg747_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg200_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg678_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1159_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1152_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1125_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1131_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1153_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1140_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1141_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1139_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1126_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product321_2_impl_1_out);

   Delay1No459_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_2_impl_1_out,
                 Y => Delay1No459_out);

Delay1No460_out_to_Product321_3_impl_parent_implementedSystem_port_0_cast <= Delay1No460_out;
Delay1No461_out_to_Product321_3_impl_parent_implementedSystem_port_1_cast <= Delay1No461_out;
   Product321_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product321_3_impl_out,
                 X => Delay1No460_out_to_Product321_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No461_out_to_Product321_3_impl_parent_implementedSystem_port_1_cast);

SharedReg862_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg862_out;
SharedReg1105_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1105_out;
SharedReg1106_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1106_out;
SharedReg1017_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1017_out;
SharedReg760_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg760_out;
SharedReg1054_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1054_out;
SharedReg990_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg990_out;
SharedReg861_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg861_out;
SharedReg683_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg683_out;
SharedReg1056_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1056_out;
SharedReg759_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg759_out;
SharedReg1158_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1158_out;
   MUX_Product321_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg862_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1105_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg759_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1158_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1106_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1017_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg760_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1054_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg990_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg861_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg683_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1056_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product321_3_impl_0_out);

   Delay1No460_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_3_impl_0_out,
                 Y => Delay1No460_out);

SharedReg1159_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1159_out;
SharedReg452_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg452_out;
SharedReg51_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg51_out;
SharedReg1152_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1152_out;
SharedReg1125_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1125_out;
SharedReg1131_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1131_out;
SharedReg1153_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1153_out;
SharedReg1140_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1140_out;
SharedReg1141_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1141_out;
SharedReg1139_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1139_out;
SharedReg1126_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1126_out;
SharedReg861_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg861_out;
   MUX_Product321_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1159_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg452_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1126_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg861_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg51_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1152_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1125_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1131_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1153_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1140_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1141_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1139_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product321_3_impl_1_out);

   Delay1No461_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_3_impl_1_out,
                 Y => Delay1No461_out);

Delay1No462_out_to_Product321_4_impl_parent_implementedSystem_port_0_cast <= Delay1No462_out;
Delay1No463_out_to_Product321_4_impl_parent_implementedSystem_port_1_cast <= Delay1No463_out;
   Product321_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product321_4_impl_out,
                 X => Delay1No462_out_to_Product321_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No463_out_to_Product321_4_impl_parent_implementedSystem_port_1_cast);

SharedReg713_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg713_out;
SharedReg1158_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1158_out;
SharedReg690_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg690_out;
SharedReg1105_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1105_out;
SharedReg1106_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1106_out;
SharedReg993_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg993_out;
SharedReg798_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg798_out;
SharedReg795_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg795_out;
SharedReg993_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg993_out;
SharedReg865_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg865_out;
SharedReg584_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg584_out;
SharedReg798_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg798_out;
   MUX_Product321_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg713_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1158_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg584_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg798_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg690_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1105_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1106_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg993_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg798_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg795_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg993_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg865_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product321_4_impl_0_out);

   Delay1No462_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_4_impl_0_out,
                 Y => Delay1No462_out);

SharedReg1126_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1126_out;
SharedReg689_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg689_out;
SharedReg1159_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1159_out;
SharedReg707_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg707_out;
SharedReg89_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg89_out;
SharedReg1152_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1152_out;
SharedReg1125_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1125_out;
SharedReg1131_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1131_out;
SharedReg1153_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1153_out;
SharedReg1140_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1140_out;
SharedReg1141_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1141_out;
SharedReg1139_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1139_out;
   MUX_Product321_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1126_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg689_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1141_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1139_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1159_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg707_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg89_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1152_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1125_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1131_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1153_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1140_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product321_4_impl_1_out);

   Delay1No463_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_4_impl_1_out,
                 Y => Delay1No463_out);

Delay1No464_out_to_Product321_5_impl_parent_implementedSystem_port_0_cast <= Delay1No464_out;
Delay1No465_out_to_Product321_5_impl_parent_implementedSystem_port_1_cast <= Delay1No465_out;
   Product321_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product321_5_impl_out,
                 X => Delay1No464_out_to_Product321_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No465_out_to_Product321_5_impl_parent_implementedSystem_port_1_cast);

SharedReg589_out_to_MUX_Product321_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg589_out;
SharedReg1062_out_to_MUX_Product321_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1062_out;
SharedReg474_out_to_MUX_Product321_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg474_out;
SharedReg1158_out_to_MUX_Product321_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1158_out;
SharedReg590_out_to_MUX_Product321_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg590_out;
SharedReg1105_out_to_MUX_Product321_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1105_out;
SharedReg1106_out_to_MUX_Product321_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1106_out;
SharedReg1028_out_to_MUX_Product321_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1028_out;
SharedReg1062_out_to_MUX_Product321_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1062_out;
SharedReg770_out_to_MUX_Product321_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg770_out;
SharedReg997_out_to_MUX_Product321_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg997_out;
SharedReg997_out_to_MUX_Product321_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg997_out;
   MUX_Product321_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg589_out_to_MUX_Product321_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1062_out_to_MUX_Product321_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg997_out_to_MUX_Product321_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg997_out_to_MUX_Product321_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg474_out_to_MUX_Product321_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1158_out_to_MUX_Product321_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg590_out_to_MUX_Product321_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1105_out_to_MUX_Product321_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1106_out_to_MUX_Product321_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1028_out_to_MUX_Product321_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1062_out_to_MUX_Product321_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg770_out_to_MUX_Product321_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product321_5_impl_0_out);

   Delay1No464_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_5_impl_0_out,
                 Y => Delay1No464_out);

SharedReg1141_out_to_MUX_Product321_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1141_out;
SharedReg1139_out_to_MUX_Product321_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1139_out;
SharedReg1126_out_to_MUX_Product321_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1126_out;
SharedReg589_out_to_MUX_Product321_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg589_out;
SharedReg1159_out_to_MUX_Product321_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1159_out;
SharedReg766_out_to_MUX_Product321_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg766_out;
SharedReg227_out_to_MUX_Product321_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg227_out;
SharedReg1152_out_to_MUX_Product321_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1152_out;
SharedReg1125_out_to_MUX_Product321_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1125_out;
SharedReg1131_out_to_MUX_Product321_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1131_out;
SharedReg1153_out_to_MUX_Product321_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1153_out;
SharedReg1140_out_to_MUX_Product321_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1140_out;
   MUX_Product321_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1141_out_to_MUX_Product321_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1139_out_to_MUX_Product321_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1153_out_to_MUX_Product321_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1140_out_to_MUX_Product321_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1126_out_to_MUX_Product321_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg589_out_to_MUX_Product321_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1159_out_to_MUX_Product321_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg766_out_to_MUX_Product321_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg227_out_to_MUX_Product321_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1152_out_to_MUX_Product321_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1125_out_to_MUX_Product321_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1131_out_to_MUX_Product321_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product321_5_impl_1_out);

   Delay1No465_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_5_impl_1_out,
                 Y => Delay1No465_out);

Delay1No466_out_to_Product321_6_impl_parent_implementedSystem_port_0_cast <= Delay1No466_out;
Delay1No467_out_to_Product321_6_impl_parent_implementedSystem_port_1_cast <= Delay1No467_out;
   Product321_6_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product321_6_impl_out,
                 X => Delay1No466_out_to_Product321_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No467_out_to_Product321_6_impl_parent_implementedSystem_port_1_cast);

SharedReg1001_out_to_MUX_Product321_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1001_out;
SharedReg871_out_to_MUX_Product321_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg871_out;
SharedReg1091_out_to_MUX_Product321_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1091_out;
SharedReg1089_out_to_MUX_Product321_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1089_out;
SharedReg1158_out_to_MUX_Product321_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1158_out;
SharedReg872_out_to_MUX_Product321_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg872_out;
SharedReg1105_out_to_MUX_Product321_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1105_out;
SharedReg1106_out_to_MUX_Product321_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1106_out;
SharedReg1075_out_to_MUX_Product321_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1075_out;
SharedReg1102_out_to_MUX_Product321_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1102_out;
SharedReg1088_out_to_MUX_Product321_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1088_out;
SharedReg1066_out_to_MUX_Product321_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1066_out;
   MUX_Product321_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1001_out_to_MUX_Product321_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg871_out_to_MUX_Product321_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1088_out_to_MUX_Product321_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1066_out_to_MUX_Product321_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1091_out_to_MUX_Product321_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1089_out_to_MUX_Product321_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1158_out_to_MUX_Product321_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg872_out_to_MUX_Product321_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1105_out_to_MUX_Product321_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1106_out_to_MUX_Product321_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1075_out_to_MUX_Product321_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1102_out_to_MUX_Product321_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product321_6_impl_0_out);

   Delay1No466_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_6_impl_0_out,
                 Y => Delay1No466_out);

SharedReg1140_out_to_MUX_Product321_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1140_out;
SharedReg1141_out_to_MUX_Product321_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1141_out;
SharedReg1139_out_to_MUX_Product321_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1139_out;
SharedReg1126_out_to_MUX_Product321_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1126_out;
SharedReg871_out_to_MUX_Product321_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg871_out;
SharedReg1159_out_to_MUX_Product321_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1159_out;
SharedReg475_out_to_MUX_Product321_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg475_out;
SharedReg391_out_to_MUX_Product321_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg391_out;
SharedReg1152_out_to_MUX_Product321_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1152_out;
SharedReg1125_out_to_MUX_Product321_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1125_out;
SharedReg1131_out_to_MUX_Product321_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1131_out;
SharedReg1153_out_to_MUX_Product321_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1153_out;
   MUX_Product321_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1140_out_to_MUX_Product321_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1141_out_to_MUX_Product321_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1131_out_to_MUX_Product321_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1153_out_to_MUX_Product321_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1139_out_to_MUX_Product321_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1126_out_to_MUX_Product321_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg871_out_to_MUX_Product321_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1159_out_to_MUX_Product321_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg475_out_to_MUX_Product321_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg391_out_to_MUX_Product321_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1152_out_to_MUX_Product321_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1125_out_to_MUX_Product321_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Product321_6_impl_1_out);

   Delay1No467_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_6_impl_1_out,
                 Y => Delay1No467_out);

Delay1No468_out_to_Subtract23_0_impl_parent_implementedSystem_port_0_cast <= Delay1No468_out;
Delay1No469_out_to_Subtract23_0_impl_parent_implementedSystem_port_1_cast <= Delay1No469_out;
   Subtract23_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract23_0_impl_out,
                 X => Delay1No468_out_to_Subtract23_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No469_out_to_Subtract23_0_impl_parent_implementedSystem_port_1_cast);

SharedReg366_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg366_out;
SharedReg4_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg7_out;
SharedReg884_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg884_out;
SharedReg530_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg530_out;
SharedReg1004_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1004_out;
SharedReg1039_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1039_out;
SharedReg1073_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1073_out;
SharedReg330_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg330_out;
SharedReg202_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg202_out;
SharedReg250_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg250_out;
Delay4No168_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_12_cast <= Delay4No168_out;
   MUX_Subtract23_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg366_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg4_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg250_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay4No168_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg7_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg884_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg530_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1004_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1039_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1073_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg330_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg202_out_to_MUX_Subtract23_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract23_0_impl_0_out);

   Delay1No468_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract23_0_impl_0_out,
                 Y => Delay1No468_out);

SharedReg371_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg371_out;
SharedReg20_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg20_out;
SharedReg23_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg23_out;
SharedReg961_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg961_out;
SharedReg625_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg625_out;
SharedReg564_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg564_out;
SharedReg670_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg670_out;
SharedReg430_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg430_out;
SharedReg363_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg363_out;
SharedReg327_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg327_out;
SharedReg363_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg363_out;
SharedReg824_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg824_out;
   MUX_Subtract23_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg371_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg20_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg363_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg824_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg23_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg961_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg625_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg564_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg670_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg430_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg363_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg327_out_to_MUX_Subtract23_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract23_0_impl_1_out);

   Delay1No469_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract23_0_impl_1_out,
                 Y => Delay1No469_out);

Delay1No470_out_to_Subtract23_1_impl_parent_implementedSystem_port_0_cast <= Delay1No470_out;
Delay1No471_out_to_Subtract23_1_impl_parent_implementedSystem_port_1_cast <= Delay1No471_out;
   Subtract23_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract23_1_impl_out,
                 X => Delay1No470_out_to_Subtract23_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No471_out_to_Subtract23_1_impl_parent_implementedSystem_port_1_cast);

SharedReg1008_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1008_out;
Delay4No169_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_2_cast <= Delay4No169_out;
SharedReg168_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg168_out;
SharedReg4_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg7_out;
SharedReg608_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg608_out;
SharedReg649_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg649_out;
SharedReg373_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg373_out;
SharedReg337_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg337_out;
SharedReg166_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg166_out;
SharedReg373_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg373_out;
SharedReg854_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg854_out;
   MUX_Subtract23_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1008_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay4No169_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg373_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg854_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg168_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg4_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg7_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg608_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg649_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg373_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg337_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg166_out_to_MUX_Subtract23_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract23_1_impl_0_out);

   Delay1No470_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract23_1_impl_0_out,
                 Y => Delay1No470_out);

Delay12No15_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_1_cast <= Delay12No15_out;
SharedReg828_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg828_out;
SharedReg380_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg380_out;
SharedReg20_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg20_out;
SharedReg23_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg23_out;
SharedReg890_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg890_out;
SharedReg826_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg826_out;
SharedReg335_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg335_out;
SharedReg379_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg379_out;
SharedReg335_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg335_out;
SharedReg164_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg164_out;
SharedReg781_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg781_out;
   MUX_Subtract23_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay12No15_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg828_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg164_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg781_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg380_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg20_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg23_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg890_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg826_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg335_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg379_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg335_out_to_MUX_Subtract23_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract23_1_impl_1_out);

   Delay1No471_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract23_1_impl_1_out,
                 Y => Delay1No471_out);

Delay1No472_out_to_Subtract23_2_impl_parent_implementedSystem_port_0_cast <= Delay1No472_out;
Delay1No473_out_to_Subtract23_2_impl_parent_implementedSystem_port_1_cast <= Delay1No473_out;
   Subtract23_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract23_2_impl_out,
                 X => Delay1No472_out_to_Subtract23_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No473_out_to_Subtract23_2_impl_parent_implementedSystem_port_1_cast);

SharedReg681_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg681_out;
SharedReg678_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg678_out;
SharedReg987_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg987_out;
Delay4No170_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_4_cast <= Delay4No170_out;
SharedReg201_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg201_out;
SharedReg5_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg5_out;
SharedReg8_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg8_out;
SharedReg893_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg893_out;
SharedReg402_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg402_out;
SharedReg445_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg445_out;
SharedReg651_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg651_out;
SharedReg76_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg76_out;
   MUX_Subtract23_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg681_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg678_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg651_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg76_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg987_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay4No170_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg201_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg5_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg8_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg893_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg402_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg445_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract23_2_impl_0_out);

   Delay1No472_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract23_2_impl_0_out,
                 Y => Delay1No472_out);

SharedReg783_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg783_out;
SharedReg788_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg788_out;
Delay12No16_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_3_cast <= Delay12No16_out;
SharedReg832_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg832_out;
SharedReg349_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg349_out;
SharedReg21_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg21_out;
SharedReg24_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg24_out;
Delay5No44_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_8_cast <= Delay5No44_out;
SharedReg510_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg510_out;
SharedReg859_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg859_out;
SharedReg829_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg829_out;
SharedReg170_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg170_out;
   MUX_Subtract23_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg783_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg788_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg829_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg170_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => Delay12No16_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg832_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg349_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg21_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg24_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay5No44_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg510_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg859_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract23_2_impl_1_out);

   Delay1No473_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract23_2_impl_1_out,
                 Y => Delay1No473_out);

Delay1No474_out_to_Subtract23_3_impl_parent_implementedSystem_port_0_cast <= Delay1No474_out;
Delay1No475_out_to_Subtract23_3_impl_parent_implementedSystem_port_1_cast <= Delay1No475_out;
   Subtract23_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract23_3_impl_out,
                 X => Delay1No474_out_to_Subtract23_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No475_out_to_Subtract23_3_impl_parent_implementedSystem_port_1_cast);

SharedReg47_out_to_MUX_Subtract23_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg47_out;
SharedReg351_out_to_MUX_Subtract23_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg351_out;
SharedReg683_out_to_MUX_Subtract23_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg683_out;
SharedReg140_out_to_MUX_Subtract23_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg140_out;
Delay4No171_out_to_MUX_Subtract23_3_impl_0_parent_implementedSystem_port_5_cast <= Delay4No171_out;
SharedReg180_out_to_MUX_Subtract23_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg180_out;
SharedReg4_out_to_MUX_Subtract23_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg4_out;
SharedReg8_out_to_MUX_Subtract23_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg8_out;
SharedReg614_out_to_MUX_Subtract23_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg614_out;
SharedReg405_out_to_MUX_Subtract23_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg405_out;
SharedReg451_out_to_MUX_Subtract23_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg451_out;
SharedReg654_out_to_MUX_Subtract23_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg654_out;
   MUX_Subtract23_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg47_out_to_MUX_Subtract23_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg351_out_to_MUX_Subtract23_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg451_out_to_MUX_Subtract23_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg654_out_to_MUX_Subtract23_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg683_out_to_MUX_Subtract23_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg140_out_to_MUX_Subtract23_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay4No171_out_to_MUX_Subtract23_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg180_out_to_MUX_Subtract23_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg4_out_to_MUX_Subtract23_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg8_out_to_MUX_Subtract23_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg614_out_to_MUX_Subtract23_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg405_out_to_MUX_Subtract23_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract23_3_impl_0_out);

   Delay1No474_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract23_3_impl_0_out,
                 Y => Delay1No474_out);

SharedReg191_out_to_MUX_Subtract23_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg191_out;
SharedReg175_out_to_MUX_Subtract23_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg175_out;
SharedReg881_out_to_MUX_Subtract23_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg881_out;
SharedReg350_out_to_MUX_Subtract23_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg350_out;
SharedReg836_out_to_MUX_Subtract23_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg836_out;
SharedReg197_out_to_MUX_Subtract23_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg197_out;
SharedReg20_out_to_MUX_Subtract23_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg20_out;
SharedReg24_out_to_MUX_Subtract23_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg24_out;
SharedReg898_out_to_MUX_Subtract23_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg898_out;
SharedReg514_out_to_MUX_Subtract23_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg514_out;
SharedReg862_out_to_MUX_Subtract23_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg862_out;
SharedReg833_out_to_MUX_Subtract23_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg833_out;
   MUX_Subtract23_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg191_out_to_MUX_Subtract23_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg175_out_to_MUX_Subtract23_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg862_out_to_MUX_Subtract23_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg833_out_to_MUX_Subtract23_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg881_out_to_MUX_Subtract23_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg350_out_to_MUX_Subtract23_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg836_out_to_MUX_Subtract23_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg197_out_to_MUX_Subtract23_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg20_out_to_MUX_Subtract23_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg24_out_to_MUX_Subtract23_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg898_out_to_MUX_Subtract23_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg514_out_to_MUX_Subtract23_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract23_3_impl_1_out);

   Delay1No475_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract23_3_impl_1_out,
                 Y => Delay1No475_out);

Delay1No476_out_to_Subtract23_4_impl_parent_implementedSystem_port_0_cast <= Delay1No476_out;
Delay1No477_out_to_Subtract23_4_impl_parent_implementedSystem_port_1_cast <= Delay1No477_out;
   Subtract23_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract23_4_impl_out,
                 X => Delay1No476_out_to_Subtract23_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No477_out_to_Subtract23_4_impl_parent_implementedSystem_port_1_cast);

SharedReg272_out_to_MUX_Subtract23_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg272_out;
SharedReg657_out_to_MUX_Subtract23_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg657_out;
SharedReg84_out_to_MUX_Subtract23_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg84_out;
SharedReg309_out_to_MUX_Subtract23_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg309_out;
SharedReg584_out_to_MUX_Subtract23_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg584_out;
SharedReg866_out_to_MUX_Subtract23_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg866_out;
Delay4No172_out_to_MUX_Subtract23_4_impl_0_parent_implementedSystem_port_7_cast <= Delay4No172_out;
SharedReg972_out_to_MUX_Subtract23_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg972_out;
SharedReg5_out_to_MUX_Subtract23_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg5_out;
SharedReg9_out_to_MUX_Subtract23_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg9_out;
SharedReg761_out_to_MUX_Subtract23_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg761_out;
SharedReg900_out_to_MUX_Subtract23_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg900_out;
   MUX_Subtract23_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg272_out_to_MUX_Subtract23_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg657_out_to_MUX_Subtract23_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg761_out_to_MUX_Subtract23_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg900_out_to_MUX_Subtract23_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg84_out_to_MUX_Subtract23_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg309_out_to_MUX_Subtract23_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg584_out_to_MUX_Subtract23_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg866_out_to_MUX_Subtract23_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay4No172_out_to_MUX_Subtract23_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg972_out_to_MUX_Subtract23_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg5_out_to_MUX_Subtract23_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg9_out_to_MUX_Subtract23_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract23_4_impl_0_out);

   Delay1No476_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract23_4_impl_0_out,
                 Y => Delay1No476_out);

SharedReg207_out_to_MUX_Subtract23_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg207_out;
SharedReg837_out_to_MUX_Subtract23_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg837_out;
SharedReg278_out_to_MUX_Subtract23_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg278_out;
SharedReg278_out_to_MUX_Subtract23_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg278_out;
SharedReg762_out_to_MUX_Subtract23_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg762_out;
Delay12No18_out_to_MUX_Subtract23_4_impl_1_parent_implementedSystem_port_6_cast <= Delay12No18_out;
SharedReg840_out_to_MUX_Subtract23_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg840_out;
SharedReg929_out_to_MUX_Subtract23_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg929_out;
SharedReg21_out_to_MUX_Subtract23_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg21_out;
SharedReg25_out_to_MUX_Subtract23_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg25_out;
SharedReg707_out_to_MUX_Subtract23_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg707_out;
SharedReg973_out_to_MUX_Subtract23_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg973_out;
   MUX_Subtract23_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg207_out_to_MUX_Subtract23_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg837_out_to_MUX_Subtract23_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg707_out_to_MUX_Subtract23_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg973_out_to_MUX_Subtract23_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg278_out_to_MUX_Subtract23_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg278_out_to_MUX_Subtract23_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg762_out_to_MUX_Subtract23_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay12No18_out_to_MUX_Subtract23_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg840_out_to_MUX_Subtract23_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg929_out_to_MUX_Subtract23_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg21_out_to_MUX_Subtract23_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg25_out_to_MUX_Subtract23_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract23_4_impl_1_out);

   Delay1No477_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract23_4_impl_1_out,
                 Y => Delay1No477_out);

Delay1No478_out_to_Subtract23_5_impl_parent_implementedSystem_port_0_cast <= Delay1No478_out;
Delay1No479_out_to_Subtract23_5_impl_parent_implementedSystem_port_1_cast <= Delay1No479_out;
   Subtract23_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract23_5_impl_out,
                 X => Delay1No478_out_to_Subtract23_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No479_out_to_Subtract23_5_impl_parent_implementedSystem_port_1_cast);

SharedReg769_out_to_MUX_Subtract23_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg769_out;
SharedReg411_out_to_MUX_Subtract23_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg411_out;
SharedReg712_out_to_MUX_Subtract23_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg712_out;
SharedReg315_out_to_MUX_Subtract23_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg315_out;
SharedReg63_out_to_MUX_Subtract23_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg63_out;
SharedReg291_out_to_MUX_Subtract23_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg291_out;
SharedReg182_out_to_MUX_Subtract23_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg182_out;
SharedReg998_out_to_MUX_Subtract23_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg998_out;
Delay4No173_out_to_MUX_Subtract23_5_impl_0_parent_implementedSystem_port_9_cast <= Delay4No173_out;
SharedReg975_out_to_MUX_Subtract23_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg975_out;
SharedReg6_out_to_MUX_Subtract23_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg6_out;
SharedReg9_out_to_MUX_Subtract23_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg9_out;
   MUX_Subtract23_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg769_out_to_MUX_Subtract23_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg411_out_to_MUX_Subtract23_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg6_out_to_MUX_Subtract23_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg9_out_to_MUX_Subtract23_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg712_out_to_MUX_Subtract23_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg315_out_to_MUX_Subtract23_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg63_out_to_MUX_Subtract23_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg291_out_to_MUX_Subtract23_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg182_out_to_MUX_Subtract23_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg998_out_to_MUX_Subtract23_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay4No173_out_to_MUX_Subtract23_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg975_out_to_MUX_Subtract23_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract23_5_impl_0_out);

   Delay1No478_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract23_5_impl_0_out,
                 Y => Delay1No478_out);

SharedReg714_out_to_MUX_Subtract23_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg714_out;
SharedReg522_out_to_MUX_Subtract23_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg522_out;
SharedReg869_out_to_MUX_Subtract23_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg869_out;
SharedReg232_out_to_MUX_Subtract23_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg232_out;
SharedReg286_out_to_MUX_Subtract23_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg286_out;
SharedReg313_out_to_MUX_Subtract23_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg313_out;
SharedReg287_out_to_MUX_Subtract23_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg287_out;
Delay12No19_out_to_MUX_Subtract23_5_impl_1_parent_implementedSystem_port_8_cast <= Delay12No19_out;
SharedReg844_out_to_MUX_Subtract23_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg844_out;
SharedReg933_out_to_MUX_Subtract23_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg933_out;
SharedReg22_out_to_MUX_Subtract23_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Subtract23_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg25_out;
   MUX_Subtract23_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg714_out_to_MUX_Subtract23_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg522_out_to_MUX_Subtract23_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg22_out_to_MUX_Subtract23_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg25_out_to_MUX_Subtract23_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg869_out_to_MUX_Subtract23_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg232_out_to_MUX_Subtract23_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg286_out_to_MUX_Subtract23_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg313_out_to_MUX_Subtract23_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg287_out_to_MUX_Subtract23_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay12No19_out_to_MUX_Subtract23_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg844_out_to_MUX_Subtract23_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg933_out_to_MUX_Subtract23_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract23_5_impl_1_out);

   Delay1No479_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract23_5_impl_1_out,
                 Y => Delay1No479_out);

Delay1No480_out_to_Subtract23_6_impl_parent_implementedSystem_port_0_cast <= Delay1No480_out;
Delay1No481_out_to_Subtract23_6_impl_parent_implementedSystem_port_1_cast <= Delay1No481_out;
   Subtract23_6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract23_6_impl_out,
                 X => Delay1No480_out_to_Subtract23_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No481_out_to_Subtract23_6_impl_parent_implementedSystem_port_1_cast);

SharedReg8_out_to_MUX_Subtract23_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg8_out;
SharedReg908_out_to_MUX_Subtract23_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg908_out;
SharedReg664_out_to_MUX_Subtract23_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg664_out;
SharedReg1033_out_to_MUX_Subtract23_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1033_out;
SharedReg1068_out_to_MUX_Subtract23_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1068_out;
SharedReg1078_out_to_MUX_Subtract23_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1078_out;
SharedReg599_out_to_MUX_Subtract23_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg599_out;
SharedReg153_out_to_MUX_Subtract23_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg153_out;
SharedReg700_out_to_MUX_Subtract23_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg700_out;
Delay4No174_out_to_MUX_Subtract23_6_impl_0_parent_implementedSystem_port_10_cast <= Delay4No174_out;
SharedReg386_out_to_MUX_Subtract23_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg386_out;
SharedReg4_out_to_MUX_Subtract23_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg4_out;
   MUX_Subtract23_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg8_out_to_MUX_Subtract23_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg908_out_to_MUX_Subtract23_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg386_out_to_MUX_Subtract23_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg4_out_to_MUX_Subtract23_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg664_out_to_MUX_Subtract23_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1033_out_to_MUX_Subtract23_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1068_out_to_MUX_Subtract23_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1078_out_to_MUX_Subtract23_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg599_out_to_MUX_Subtract23_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg153_out_to_MUX_Subtract23_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg700_out_to_MUX_Subtract23_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay4No174_out_to_MUX_Subtract23_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract23_6_impl_0_out);

   Delay1No480_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract23_6_impl_0_out,
                 Y => Delay1No480_out);

SharedReg24_out_to_MUX_Subtract23_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg24_out;
SharedReg979_out_to_MUX_Subtract23_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg979_out;
SharedReg846_out_to_MUX_Subtract23_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg846_out;
SharedReg595_out_to_MUX_Subtract23_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg595_out;
SharedReg704_out_to_MUX_Subtract23_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg704_out;
SharedReg770_out_to_MUX_Subtract23_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg770_out;
SharedReg1066_out_to_MUX_Subtract23_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1066_out;
SharedReg356_out_to_MUX_Subtract23_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg356_out;
SharedReg871_out_to_MUX_Subtract23_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg871_out;
SharedReg848_out_to_MUX_Subtract23_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg848_out;
SharedReg394_out_to_MUX_Subtract23_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg394_out;
SharedReg20_out_to_MUX_Subtract23_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg20_out;
   MUX_Subtract23_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg24_out_to_MUX_Subtract23_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg979_out_to_MUX_Subtract23_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg394_out_to_MUX_Subtract23_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg20_out_to_MUX_Subtract23_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg846_out_to_MUX_Subtract23_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg595_out_to_MUX_Subtract23_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg704_out_to_MUX_Subtract23_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg770_out_to_MUX_Subtract23_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1066_out_to_MUX_Subtract23_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg356_out_to_MUX_Subtract23_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg871_out_to_MUX_Subtract23_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg848_out_to_MUX_Subtract23_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract23_6_impl_1_out);

   Delay1No481_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract23_6_impl_1_out,
                 Y => Delay1No481_out);

Delay1No482_out_to_Subtract30_0_impl_parent_implementedSystem_port_0_cast <= Delay1No482_out;
Delay1No483_out_to_Subtract30_0_impl_parent_implementedSystem_port_1_cast <= Delay1No483_out;
   Subtract30_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract30_0_impl_out,
                 X => Delay1No482_out_to_Subtract30_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No483_out_to_Subtract30_0_impl_parent_implementedSystem_port_1_cast);

SharedReg960_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg960_out;
SharedReg5_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg5_out;
SharedReg8_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg8_out;
SharedReg605_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg605_out;
SharedReg646_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg646_out;
SharedReg327_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg327_out;
SharedReg298_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg298_out;
SharedReg365_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg365_out;
SharedReg327_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg327_out;
SharedReg981_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg981_out;
SharedReg1038_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1038_out;
SharedReg531_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg531_out;
   MUX_Subtract30_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg960_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg5_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1038_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg531_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg8_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg605_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg646_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg327_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg298_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg365_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg327_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg981_out_to_MUX_Subtract30_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract30_0_impl_0_out);

   Delay1No482_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract30_0_impl_0_out,
                 Y => Delay1No482_out);

SharedReg913_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg913_out;
SharedReg21_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg21_out;
SharedReg24_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg24_out;
SharedReg886_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg886_out;
SharedReg822_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg822_out;
SharedReg297_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg297_out;
SharedReg370_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg370_out;
SharedReg297_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg297_out;
SharedReg158_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg158_out;
SharedReg436_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg436_out;
Delay12No14_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_11_cast <= Delay12No14_out;
SharedReg626_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg626_out;
   MUX_Subtract30_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg913_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg21_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay12No14_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg626_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg24_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg886_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg822_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg297_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg370_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg297_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg158_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg436_out_to_MUX_Subtract30_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract30_0_impl_1_out);

   Delay1No483_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract30_0_impl_1_out,
                 Y => Delay1No483_out);

Delay1No484_out_to_Subtract30_1_impl_parent_implementedSystem_port_0_cast <= Delay1No484_out;
Delay1No485_out_to_Subtract30_1_impl_parent_implementedSystem_port_1_cast <= Delay1No485_out;
   Subtract30_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract30_1_impl_out,
                 X => Delay1No484_out_to_Subtract30_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No485_out_to_Subtract30_1_impl_parent_implementedSystem_port_1_cast);

SharedReg373_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg373_out;
SharedReg534_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg534_out;
SharedReg963_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg963_out;
SharedReg5_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg5_out;
SharedReg8_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg8_out;
SharedReg889_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg889_out;
SharedReg399_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg399_out;
SharedReg438_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg438_out;
SharedReg648_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg648_out;
SharedReg40_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg40_out;
SharedReg675_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg675_out;
SharedReg254_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg254_out;
   MUX_Subtract30_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg373_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg534_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg675_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg254_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg963_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg5_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg8_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg889_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg399_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg438_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg648_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg40_out_to_MUX_Subtract30_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract30_1_impl_0_out);

   Delay1No484_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract30_1_impl_0_out,
                 Y => Delay1No484_out);

SharedReg340_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg340_out;
SharedReg629_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg629_out;
SharedReg917_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg917_out;
SharedReg21_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg21_out;
SharedReg24_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg24_out;
Delay5No43_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_6_cast <= Delay5No43_out;
SharedReg506_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg506_out;
SharedReg855_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg855_out;
SharedReg825_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg825_out;
SharedReg164_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg164_out;
SharedReg775_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg775_out;
SharedReg237_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg237_out;
   MUX_Subtract30_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg340_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg629_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg775_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg237_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg917_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg21_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg24_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay5No43_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg506_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg855_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg825_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg164_out_to_MUX_Subtract30_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract30_1_impl_1_out);

   Delay1No485_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract30_1_impl_1_out,
                 Y => Delay1No485_out);

Delay1No486_out_to_Subtract30_2_impl_parent_implementedSystem_port_0_cast <= Delay1No486_out;
Delay1No487_out_to_Subtract30_2_impl_parent_implementedSystem_port_1_cast <= Delay1No487_out;
   Subtract30_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract30_2_impl_out,
                 X => Delay1No486_out_to_Subtract30_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No487_out_to_Subtract30_2_impl_parent_implementedSystem_port_1_cast);

SharedReg137_out_to_MUX_Subtract30_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg137_out;
SharedReg260_out_to_MUX_Subtract30_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg260_out;
SharedReg343_out_to_MUX_Subtract30_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg343_out;
SharedReg537_out_to_MUX_Subtract30_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg537_out;
SharedReg966_out_to_MUX_Subtract30_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg966_out;
SharedReg6_out_to_MUX_Subtract30_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg6_out;
SharedReg9_out_to_MUX_Subtract30_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg9_out;
SharedReg750_out_to_MUX_Subtract30_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg750_out;
SharedReg892_out_to_MUX_Subtract30_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg892_out;
SharedReg302_out_to_MUX_Subtract30_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg302_out;
SharedReg891_out_to_MUX_Subtract30_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg891_out;
SharedReg578_out_to_MUX_Subtract30_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg578_out;
   MUX_Subtract30_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg137_out_to_MUX_Subtract30_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg260_out_to_MUX_Subtract30_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg891_out_to_MUX_Subtract30_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg578_out_to_MUX_Subtract30_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg343_out_to_MUX_Subtract30_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg537_out_to_MUX_Subtract30_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg966_out_to_MUX_Subtract30_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg6_out_to_MUX_Subtract30_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg9_out_to_MUX_Subtract30_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg750_out_to_MUX_Subtract30_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg892_out_to_MUX_Subtract30_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg302_out_to_MUX_Subtract30_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract30_2_impl_0_out);

   Delay1No486_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract30_2_impl_0_out,
                 Y => Delay1No486_out);

SharedReg134_out_to_MUX_Subtract30_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg134_out;
SharedReg242_out_to_MUX_Subtract30_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg242_out;
SharedReg306_out_to_MUX_Subtract30_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg306_out;
SharedReg632_out_to_MUX_Subtract30_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg632_out;
SharedReg921_out_to_MUX_Subtract30_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg921_out;
SharedReg22_out_to_MUX_Subtract30_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Subtract30_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg25_out;
SharedReg785_out_to_MUX_Subtract30_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg785_out;
SharedReg967_out_to_MUX_Subtract30_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg967_out;
SharedReg240_out_to_MUX_Subtract30_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg240_out;
SharedReg966_out_to_MUX_Subtract30_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg966_out;
SharedReg576_out_to_MUX_Subtract30_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg576_out;
   MUX_Subtract30_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg134_out_to_MUX_Subtract30_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg242_out_to_MUX_Subtract30_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg966_out_to_MUX_Subtract30_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg576_out_to_MUX_Subtract30_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg306_out_to_MUX_Subtract30_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg632_out_to_MUX_Subtract30_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg921_out_to_MUX_Subtract30_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg22_out_to_MUX_Subtract30_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg25_out_to_MUX_Subtract30_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg785_out_to_MUX_Subtract30_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg967_out_to_MUX_Subtract30_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg240_out_to_MUX_Subtract30_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract30_2_impl_1_out);

   Delay1No487_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract30_2_impl_1_out,
                 Y => Delay1No487_out);

Delay1No488_out_to_Subtract30_3_impl_parent_implementedSystem_port_0_cast <= Delay1No488_out;
Delay1No489_out_to_Subtract30_3_impl_parent_implementedSystem_port_1_cast <= Delay1No489_out;
   Subtract30_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract30_3_impl_out,
                 X => Delay1No488_out_to_Subtract30_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No489_out_to_Subtract30_3_impl_parent_implementedSystem_port_1_cast);

SharedReg582_out_to_MUX_Subtract30_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg582_out;
SharedReg686_out_to_MUX_Subtract30_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg686_out;
SharedReg244_out_to_MUX_Subtract30_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg244_out;
SharedReg991_out_to_MUX_Subtract30_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg991_out;
SharedReg540_out_to_MUX_Subtract30_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg540_out;
SharedReg969_out_to_MUX_Subtract30_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg969_out;
SharedReg5_out_to_MUX_Subtract30_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg5_out;
SharedReg9_out_to_MUX_Subtract30_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg9_out;
SharedReg897_out_to_MUX_Subtract30_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg897_out;
SharedReg896_out_to_MUX_Subtract30_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg896_out;
SharedReg266_out_to_MUX_Subtract30_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg266_out;
SharedReg895_out_to_MUX_Subtract30_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg895_out;
   MUX_Subtract30_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg582_out_to_MUX_Subtract30_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg686_out_to_MUX_Subtract30_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg266_out_to_MUX_Subtract30_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg895_out_to_MUX_Subtract30_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg244_out_to_MUX_Subtract30_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg991_out_to_MUX_Subtract30_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg540_out_to_MUX_Subtract30_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg969_out_to_MUX_Subtract30_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg5_out_to_MUX_Subtract30_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg9_out_to_MUX_Subtract30_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg897_out_to_MUX_Subtract30_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg896_out_to_MUX_Subtract30_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract30_3_impl_0_out);

   Delay1No488_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract30_3_impl_0_out,
                 Y => Delay1No488_out);

SharedReg580_out_to_MUX_Subtract30_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg580_out;
SharedReg753_out_to_MUX_Subtract30_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg753_out;
SharedReg143_out_to_MUX_Subtract30_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg143_out;
Delay12No17_out_to_MUX_Subtract30_3_impl_1_parent_implementedSystem_port_4_cast <= Delay12No17_out;
SharedReg635_out_to_MUX_Subtract30_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg635_out;
SharedReg925_out_to_MUX_Subtract30_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg925_out;
SharedReg21_out_to_MUX_Subtract30_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg21_out;
SharedReg25_out_to_MUX_Subtract30_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg25_out;
Delay5No45_out_to_MUX_Subtract30_3_impl_1_parent_implementedSystem_port_9_cast <= Delay5No45_out;
SharedReg970_out_to_MUX_Subtract30_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg970_out;
SharedReg140_out_to_MUX_Subtract30_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg140_out;
SharedReg969_out_to_MUX_Subtract30_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg969_out;
   MUX_Subtract30_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg580_out_to_MUX_Subtract30_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg753_out_to_MUX_Subtract30_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg140_out_to_MUX_Subtract30_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg969_out_to_MUX_Subtract30_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg143_out_to_MUX_Subtract30_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay12No17_out_to_MUX_Subtract30_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg635_out_to_MUX_Subtract30_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg925_out_to_MUX_Subtract30_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg21_out_to_MUX_Subtract30_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg25_out_to_MUX_Subtract30_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay5No45_out_to_MUX_Subtract30_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg970_out_to_MUX_Subtract30_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract30_3_impl_1_out);

   Delay1No489_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract30_3_impl_1_out,
                 Y => Delay1No489_out);

Delay1No490_out_to_Subtract30_4_impl_parent_implementedSystem_port_0_cast <= Delay1No490_out;
Delay1No491_out_to_Subtract30_4_impl_parent_implementedSystem_port_1_cast <= Delay1No491_out;
   Subtract30_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract30_4_impl_out,
                 X => Delay1No490_out_to_Subtract30_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No491_out_to_Subtract30_4_impl_parent_implementedSystem_port_1_cast);

SharedReg709_out_to_MUX_Subtract30_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg709_out;
SharedReg899_out_to_MUX_Subtract30_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg899_out;
SharedReg586_out_to_MUX_Subtract30_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg586_out;
SharedReg692_out_to_MUX_Subtract30_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg692_out;
SharedReg206_out_to_MUX_Subtract30_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg206_out;
SharedReg309_out_to_MUX_Subtract30_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg309_out;
SharedReg543_out_to_MUX_Subtract30_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg543_out;
SharedReg587_out_to_MUX_Subtract30_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg587_out;
SharedReg6_out_to_MUX_Subtract30_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg6_out;
SharedReg11_out_to_MUX_Subtract30_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg11_out;
SharedReg85_out_to_MUX_Subtract30_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg85_out;
SharedReg794_out_to_MUX_Subtract30_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg794_out;
   MUX_Subtract30_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg709_out_to_MUX_Subtract30_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg899_out_to_MUX_Subtract30_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg85_out_to_MUX_Subtract30_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg794_out_to_MUX_Subtract30_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg586_out_to_MUX_Subtract30_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg692_out_to_MUX_Subtract30_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg206_out_to_MUX_Subtract30_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg309_out_to_MUX_Subtract30_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg543_out_to_MUX_Subtract30_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg587_out_to_MUX_Subtract30_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg6_out_to_MUX_Subtract30_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg11_out_to_MUX_Subtract30_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract30_4_impl_0_out);

   Delay1No490_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract30_4_impl_0_out,
                 Y => Delay1No490_out);

SharedReg994_out_to_MUX_Subtract30_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg994_out;
SharedReg972_out_to_MUX_Subtract30_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg972_out;
SharedReg458_out_to_MUX_Subtract30_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg458_out;
SharedReg790_out_to_MUX_Subtract30_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg790_out;
SharedReg211_out_to_MUX_Subtract30_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg211_out;
SharedReg311_out_to_MUX_Subtract30_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg311_out;
SharedReg638_out_to_MUX_Subtract30_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg638_out;
SharedReg763_out_to_MUX_Subtract30_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg763_out;
SharedReg22_out_to_MUX_Subtract30_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg22_out;
SharedReg27_out_to_MUX_Subtract30_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg27_out;
SharedReg310_out_to_MUX_Subtract30_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg310_out;
SharedReg707_out_to_MUX_Subtract30_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg707_out;
   MUX_Subtract30_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg994_out_to_MUX_Subtract30_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg972_out_to_MUX_Subtract30_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg310_out_to_MUX_Subtract30_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg707_out_to_MUX_Subtract30_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg458_out_to_MUX_Subtract30_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg790_out_to_MUX_Subtract30_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg211_out_to_MUX_Subtract30_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg311_out_to_MUX_Subtract30_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg638_out_to_MUX_Subtract30_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg763_out_to_MUX_Subtract30_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg22_out_to_MUX_Subtract30_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg27_out_to_MUX_Subtract30_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract30_4_impl_1_out);

   Delay1No491_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract30_4_impl_1_out,
                 Y => Delay1No491_out);

Delay1No492_out_to_Subtract30_5_impl_parent_implementedSystem_port_0_cast <= Delay1No492_out;
Delay1No493_out_to_Subtract30_5_impl_parent_implementedSystem_port_1_cast <= Delay1No493_out;
   Subtract30_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract30_5_impl_out,
                 X => Delay1No492_out_to_Subtract30_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No493_out_to_Subtract30_5_impl_parent_implementedSystem_port_1_cast);

SharedReg122_out_to_MUX_Subtract30_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg122_out;
SharedReg904_out_to_MUX_Subtract30_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg904_out;
SharedReg286_out_to_MUX_Subtract30_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg286_out;
SharedReg660_out_to_MUX_Subtract30_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg660_out;
SharedReg121_out_to_MUX_Subtract30_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg121_out;
SharedReg697_out_to_MUX_Subtract30_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg697_out;
SharedReg694_out_to_MUX_Subtract30_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg694_out;
SharedReg314_out_to_MUX_Subtract30_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg314_out;
SharedReg546_out_to_MUX_Subtract30_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg546_out;
SharedReg592_out_to_MUX_Subtract30_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg592_out;
SharedReg10_out_to_MUX_Subtract30_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg10_out;
SharedReg11_out_to_MUX_Subtract30_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg11_out;
   MUX_Subtract30_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg122_out_to_MUX_Subtract30_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg904_out_to_MUX_Subtract30_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg10_out_to_MUX_Subtract30_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg11_out_to_MUX_Subtract30_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg286_out_to_MUX_Subtract30_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg660_out_to_MUX_Subtract30_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg121_out_to_MUX_Subtract30_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg697_out_to_MUX_Subtract30_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg694_out_to_MUX_Subtract30_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg314_out_to_MUX_Subtract30_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg546_out_to_MUX_Subtract30_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg592_out_to_MUX_Subtract30_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract30_5_impl_0_out);

   Delay1No492_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract30_5_impl_0_out,
                 Y => Delay1No492_out);

SharedReg292_out_to_MUX_Subtract30_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg292_out;
SharedReg976_out_to_MUX_Subtract30_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg976_out;
SharedReg213_out_to_MUX_Subtract30_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg213_out;
SharedReg841_out_to_MUX_Subtract30_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg841_out;
SharedReg313_out_to_MUX_Subtract30_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg313_out;
SharedReg795_out_to_MUX_Subtract30_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg795_out;
SharedReg716_out_to_MUX_Subtract30_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg716_out;
SharedReg318_out_to_MUX_Subtract30_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg318_out;
SharedReg641_out_to_MUX_Subtract30_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg641_out;
SharedReg717_out_to_MUX_Subtract30_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg717_out;
SharedReg26_out_to_MUX_Subtract30_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg26_out;
SharedReg27_out_to_MUX_Subtract30_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg27_out;
   MUX_Subtract30_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg292_out_to_MUX_Subtract30_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg976_out_to_MUX_Subtract30_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg26_out_to_MUX_Subtract30_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg27_out_to_MUX_Subtract30_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg213_out_to_MUX_Subtract30_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg841_out_to_MUX_Subtract30_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg313_out_to_MUX_Subtract30_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg795_out_to_MUX_Subtract30_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg716_out_to_MUX_Subtract30_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg318_out_to_MUX_Subtract30_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg641_out_to_MUX_Subtract30_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg717_out_to_MUX_Subtract30_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract30_5_impl_1_out);

   Delay1No493_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract30_5_impl_1_out,
                 Y => Delay1No493_out);

Delay1No494_out_to_Subtract30_6_impl_parent_implementedSystem_port_0_cast <= Delay1No494_out;
Delay1No495_out_to_Subtract30_6_impl_parent_implementedSystem_port_1_cast <= Delay1No495_out;
   Subtract30_6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract30_6_impl_out,
                 X => Delay1No494_out_to_Subtract30_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No495_out_to_Subtract30_6_impl_parent_implementedSystem_port_1_cast);

SharedReg9_out_to_MUX_Subtract30_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg9_out;
SharedReg623_out_to_MUX_Subtract30_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg623_out;
SharedReg414_out_to_MUX_Subtract30_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg414_out;
SharedReg356_out_to_MUX_Subtract30_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg356_out;
SharedReg322_out_to_MUX_Subtract30_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg322_out;
SharedReg384_out_to_MUX_Subtract30_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg384_out;
SharedReg385_out_to_MUX_Subtract30_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg385_out;
SharedReg871_out_to_MUX_Subtract30_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg871_out;
SharedReg188_out_to_MUX_Subtract30_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg188_out;
SharedReg549_out_to_MUX_Subtract30_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg549_out;
SharedReg978_out_to_MUX_Subtract30_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg978_out;
SharedReg5_out_to_MUX_Subtract30_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg5_out;
   MUX_Subtract30_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg9_out_to_MUX_Subtract30_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg623_out_to_MUX_Subtract30_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg978_out_to_MUX_Subtract30_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg5_out_to_MUX_Subtract30_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg414_out_to_MUX_Subtract30_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg356_out_to_MUX_Subtract30_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg322_out_to_MUX_Subtract30_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg384_out_to_MUX_Subtract30_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg385_out_to_MUX_Subtract30_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg871_out_to_MUX_Subtract30_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg188_out_to_MUX_Subtract30_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg549_out_to_MUX_Subtract30_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract30_6_impl_0_out);

   Delay1No494_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract30_6_impl_0_out,
                 Y => Delay1No494_out);

SharedReg25_out_to_MUX_Subtract30_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg25_out;
SharedReg910_out_to_MUX_Subtract30_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg910_out;
SharedReg526_out_to_MUX_Subtract30_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg526_out;
SharedReg320_out_to_MUX_Subtract30_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg320_out;
SharedReg388_out_to_MUX_Subtract30_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg388_out;
SharedReg218_out_to_MUX_Subtract30_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg218_out;
SharedReg381_out_to_MUX_Subtract30_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg381_out;
SharedReg478_out_to_MUX_Subtract30_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg478_out;
SharedReg381_out_to_MUX_Subtract30_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg381_out;
SharedReg644_out_to_MUX_Subtract30_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg644_out;
SharedReg937_out_to_MUX_Subtract30_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg937_out;
SharedReg21_out_to_MUX_Subtract30_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg21_out;
   MUX_Subtract30_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg25_out_to_MUX_Subtract30_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg910_out_to_MUX_Subtract30_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg937_out_to_MUX_Subtract30_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg21_out_to_MUX_Subtract30_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg526_out_to_MUX_Subtract30_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg320_out_to_MUX_Subtract30_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg388_out_to_MUX_Subtract30_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg218_out_to_MUX_Subtract30_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg381_out_to_MUX_Subtract30_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg478_out_to_MUX_Subtract30_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg381_out_to_MUX_Subtract30_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg644_out_to_MUX_Subtract30_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract30_6_impl_1_out);

   Delay1No495_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract30_6_impl_1_out,
                 Y => Delay1No495_out);

Delay1No496_out_to_Subtract32_0_impl_parent_implementedSystem_port_0_cast <= Delay1No496_out;
Delay1No497_out_to_Subtract32_0_impl_parent_implementedSystem_port_1_cast <= Delay1No497_out;
   Subtract32_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract32_0_impl_out,
                 X => Delay1No496_out_to_Subtract32_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No497_out_to_Subtract32_0_impl_parent_implementedSystem_port_1_cast);

SharedReg669_out_to_MUX_Subtract32_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg669_out;
SharedReg6_out_to_MUX_Subtract32_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg6_out;
SharedReg9_out_to_MUX_Subtract32_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg9_out;
SharedReg885_out_to_MUX_Subtract32_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg885_out;
SharedReg396_out_to_MUX_Subtract32_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg396_out;
SharedReg430_out_to_MUX_Subtract32_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg430_out;
SharedReg645_out_to_MUX_Subtract32_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg645_out;
SharedReg35_out_to_MUX_Subtract32_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg35_out;
SharedReg668_out_to_MUX_Subtract32_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg668_out;
SharedReg297_out_to_MUX_Subtract32_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg297_out;
SharedReg364_out_to_MUX_Subtract32_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg364_out;
SharedReg647_out_to_MUX_Subtract32_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg647_out;
   MUX_Subtract32_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg669_out_to_MUX_Subtract32_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg6_out_to_MUX_Subtract32_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg364_out_to_MUX_Subtract32_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg647_out_to_MUX_Subtract32_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg9_out_to_MUX_Subtract32_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg885_out_to_MUX_Subtract32_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg396_out_to_MUX_Subtract32_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg430_out_to_MUX_Subtract32_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg645_out_to_MUX_Subtract32_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg35_out_to_MUX_Subtract32_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg668_out_to_MUX_Subtract32_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg297_out_to_MUX_Subtract32_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract32_0_impl_0_out);

   Delay1No496_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract32_0_impl_0_out,
                 Y => Delay1No496_out);

SharedReg437_out_to_MUX_Subtract32_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg437_out;
SharedReg22_out_to_MUX_Subtract32_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Subtract32_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg25_out;
Delay5No42_out_to_MUX_Subtract32_0_impl_1_parent_implementedSystem_port_4_cast <= Delay5No42_out;
SharedReg502_out_to_MUX_Subtract32_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg502_out;
SharedReg850_out_to_MUX_Subtract32_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg850_out;
SharedReg821_out_to_MUX_Subtract32_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg821_out;
SharedReg363_out_to_MUX_Subtract32_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg363_out;
SharedReg430_out_to_MUX_Subtract32_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg430_out;
SharedReg252_out_to_MUX_Subtract32_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg252_out;
SharedReg333_out_to_MUX_Subtract32_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg333_out;
SharedReg823_out_to_MUX_Subtract32_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg823_out;
   MUX_Subtract32_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg437_out_to_MUX_Subtract32_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg22_out_to_MUX_Subtract32_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg333_out_to_MUX_Subtract32_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg823_out_to_MUX_Subtract32_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg25_out_to_MUX_Subtract32_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay5No42_out_to_MUX_Subtract32_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg502_out_to_MUX_Subtract32_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg850_out_to_MUX_Subtract32_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg821_out_to_MUX_Subtract32_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg363_out_to_MUX_Subtract32_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg430_out_to_MUX_Subtract32_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg252_out_to_MUX_Subtract32_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract32_0_impl_1_out);

   Delay1No497_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract32_0_impl_1_out,
                 Y => Delay1No497_out);

Delay1No498_out_to_Subtract32_1_impl_parent_implementedSystem_port_0_cast <= Delay1No498_out;
Delay1No499_out_to_Subtract32_1_impl_parent_implementedSystem_port_1_cast <= Delay1No499_out;
   Subtract32_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract32_1_impl_out,
                 X => Delay1No498_out_to_Subtract32_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No499_out_to_Subtract32_1_impl_parent_implementedSystem_port_1_cast);

SharedReg1043_out_to_MUX_Subtract32_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1043_out;
SharedReg650_out_to_MUX_Subtract32_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg650_out;
SharedReg676_out_to_MUX_Subtract32_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg676_out;
SharedReg6_out_to_MUX_Subtract32_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg6_out;
SharedReg9_out_to_MUX_Subtract32_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg9_out;
SharedReg442_out_to_MUX_Subtract32_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg442_out;
SharedReg888_out_to_MUX_Subtract32_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg888_out;
SharedReg254_out_to_MUX_Subtract32_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg254_out;
SharedReg887_out_to_MUX_Subtract32_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg887_out;
SharedReg572_out_to_MUX_Subtract32_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg572_out;
SharedReg103_out_to_MUX_Subtract32_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg103_out;
SharedReg984_out_to_MUX_Subtract32_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg984_out;
   MUX_Subtract32_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1043_out_to_MUX_Subtract32_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg650_out_to_MUX_Subtract32_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg103_out_to_MUX_Subtract32_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg984_out_to_MUX_Subtract32_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg676_out_to_MUX_Subtract32_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg6_out_to_MUX_Subtract32_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg9_out_to_MUX_Subtract32_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg442_out_to_MUX_Subtract32_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg888_out_to_MUX_Subtract32_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg254_out_to_MUX_Subtract32_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg887_out_to_MUX_Subtract32_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg572_out_to_MUX_Subtract32_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract32_1_impl_0_out);

   Delay1No498_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract32_1_impl_0_out,
                 Y => Delay1No498_out);

SharedReg1046_out_to_MUX_Subtract32_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1046_out;
SharedReg827_out_to_MUX_Subtract32_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg827_out;
SharedReg782_out_to_MUX_Subtract32_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg782_out;
SharedReg22_out_to_MUX_Subtract32_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Subtract32_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg25_out;
SharedReg777_out_to_MUX_Subtract32_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg777_out;
SharedReg964_out_to_MUX_Subtract32_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg964_out;
SharedReg131_out_to_MUX_Subtract32_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg131_out;
SharedReg963_out_to_MUX_Subtract32_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg963_out;
SharedReg672_out_to_MUX_Subtract32_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg672_out;
SharedReg130_out_to_MUX_Subtract32_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg130_out;
SharedReg443_out_to_MUX_Subtract32_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg443_out;
   MUX_Subtract32_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1046_out_to_MUX_Subtract32_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg827_out_to_MUX_Subtract32_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg130_out_to_MUX_Subtract32_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg443_out_to_MUX_Subtract32_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg782_out_to_MUX_Subtract32_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg22_out_to_MUX_Subtract32_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg25_out_to_MUX_Subtract32_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg777_out_to_MUX_Subtract32_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg964_out_to_MUX_Subtract32_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg131_out_to_MUX_Subtract32_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg963_out_to_MUX_Subtract32_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg672_out_to_MUX_Subtract32_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract32_1_impl_1_out);

   Delay1No499_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract32_1_impl_1_out,
                 Y => Delay1No499_out);

Delay1No500_out_to_Subtract32_2_impl_parent_implementedSystem_port_0_cast <= Delay1No500_out;
Delay1No501_out_to_Subtract32_2_impl_parent_implementedSystem_port_1_cast <= Delay1No501_out;
   Subtract32_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract32_2_impl_out,
                 X => Delay1No500_out_to_Subtract32_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No501_out_to_Subtract32_2_impl_parent_implementedSystem_port_1_cast);

SharedReg447_out_to_MUX_Subtract32_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg447_out;
SharedReg858_out_to_MUX_Subtract32_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg858_out;
SharedReg1013_out_to_MUX_Subtract32_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1013_out;
SharedReg653_out_to_MUX_Subtract32_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg653_out;
SharedReg682_out_to_MUX_Subtract32_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg682_out;
SharedReg10_out_to_MUX_Subtract32_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg10_out;
SharedReg11_out_to_MUX_Subtract32_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg11_out;
SharedReg109_out_to_MUX_Subtract32_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg109_out;
SharedReg787_out_to_MUX_Subtract32_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg787_out;
SharedReg448_out_to_MUX_Subtract32_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg448_out;
SharedReg305_out_to_MUX_Subtract32_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg305_out;
SharedReg108_out_to_MUX_Subtract32_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg108_out;
   MUX_Subtract32_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg447_out_to_MUX_Subtract32_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg858_out_to_MUX_Subtract32_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg305_out_to_MUX_Subtract32_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg108_out_to_MUX_Subtract32_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1013_out_to_MUX_Subtract32_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg653_out_to_MUX_Subtract32_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg682_out_to_MUX_Subtract32_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg10_out_to_MUX_Subtract32_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg11_out_to_MUX_Subtract32_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg109_out_to_MUX_Subtract32_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg787_out_to_MUX_Subtract32_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg448_out_to_MUX_Subtract32_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract32_2_impl_0_out);

   Delay1No500_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract32_2_impl_0_out,
                 Y => Delay1No500_out);

SharedReg858_out_to_MUX_Subtract32_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg858_out;
SharedReg751_out_to_MUX_Subtract32_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg751_out;
SharedReg1016_out_to_MUX_Subtract32_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1016_out;
SharedReg831_out_to_MUX_Subtract32_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg831_out;
SharedReg789_out_to_MUX_Subtract32_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg789_out;
SharedReg26_out_to_MUX_Subtract32_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg26_out;
SharedReg27_out_to_MUX_Subtract32_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg27_out;
SharedReg262_out_to_MUX_Subtract32_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg262_out;
SharedReg747_out_to_MUX_Subtract32_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg747_out;
SharedReg987_out_to_MUX_Subtract32_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg987_out;
SharedReg262_out_to_MUX_Subtract32_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg262_out;
SharedReg198_out_to_MUX_Subtract32_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg198_out;
   MUX_Subtract32_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg858_out_to_MUX_Subtract32_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg751_out_to_MUX_Subtract32_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg262_out_to_MUX_Subtract32_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg198_out_to_MUX_Subtract32_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg1016_out_to_MUX_Subtract32_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg831_out_to_MUX_Subtract32_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg789_out_to_MUX_Subtract32_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg26_out_to_MUX_Subtract32_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg27_out_to_MUX_Subtract32_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg262_out_to_MUX_Subtract32_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg747_out_to_MUX_Subtract32_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg987_out_to_MUX_Subtract32_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract32_2_impl_1_out);

   Delay1No501_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract32_2_impl_1_out,
                 Y => Delay1No501_out);

Delay1No502_out_to_Subtract32_3_impl_parent_implementedSystem_port_0_cast <= Delay1No502_out;
Delay1No503_out_to_Subtract32_3_impl_parent_implementedSystem_port_1_cast <= Delay1No503_out;
   Subtract32_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract32_3_impl_out,
                 X => Delay1No502_out_to_Subtract32_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No503_out_to_Subtract32_3_impl_parent_implementedSystem_port_1_cast);

SharedReg80_out_to_MUX_Subtract32_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg80_out;
SharedReg112_out_to_MUX_Subtract32_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg112_out;
SharedReg861_out_to_MUX_Subtract32_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg861_out;
SharedReg351_out_to_MUX_Subtract32_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg351_out;
SharedReg656_out_to_MUX_Subtract32_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg656_out;
SharedReg687_out_to_MUX_Subtract32_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg687_out;
SharedReg6_out_to_MUX_Subtract32_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg6_out;
SharedReg11_out_to_MUX_Subtract32_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg11_out;
SharedReg456_out_to_MUX_Subtract32_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg456_out;
SharedReg880_out_to_MUX_Subtract32_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg880_out;
SharedReg456_out_to_MUX_Subtract32_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg456_out;
SharedReg269_out_to_MUX_Subtract32_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg269_out;
   MUX_Subtract32_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg80_out_to_MUX_Subtract32_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg112_out_to_MUX_Subtract32_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg456_out_to_MUX_Subtract32_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg269_out_to_MUX_Subtract32_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg861_out_to_MUX_Subtract32_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg351_out_to_MUX_Subtract32_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg656_out_to_MUX_Subtract32_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg687_out_to_MUX_Subtract32_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg6_out_to_MUX_Subtract32_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg11_out_to_MUX_Subtract32_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg456_out_to_MUX_Subtract32_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg880_out_to_MUX_Subtract32_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract32_3_impl_0_out);

   Delay1No502_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract32_3_impl_0_out,
                 Y => Delay1No502_out);

SharedReg175_out_to_MUX_Subtract32_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg175_out;
SharedReg139_out_to_MUX_Subtract32_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg139_out;
SharedReg756_out_to_MUX_Subtract32_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg756_out;
SharedReg270_out_to_MUX_Subtract32_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg270_out;
SharedReg835_out_to_MUX_Subtract32_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg835_out;
SharedReg882_out_to_MUX_Subtract32_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg882_out;
SharedReg22_out_to_MUX_Subtract32_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg22_out;
SharedReg27_out_to_MUX_Subtract32_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg27_out;
SharedReg755_out_to_MUX_Subtract32_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg755_out;
SharedReg755_out_to_MUX_Subtract32_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg755_out;
SharedReg991_out_to_MUX_Subtract32_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg991_out;
SharedReg246_out_to_MUX_Subtract32_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg246_out;
   MUX_Subtract32_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg175_out_to_MUX_Subtract32_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg139_out_to_MUX_Subtract32_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg991_out_to_MUX_Subtract32_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg246_out_to_MUX_Subtract32_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg756_out_to_MUX_Subtract32_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg270_out_to_MUX_Subtract32_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg835_out_to_MUX_Subtract32_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg882_out_to_MUX_Subtract32_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg22_out_to_MUX_Subtract32_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg27_out_to_MUX_Subtract32_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg755_out_to_MUX_Subtract32_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg755_out_to_MUX_Subtract32_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract32_3_impl_1_out);

   Delay1No503_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract32_3_impl_1_out,
                 Y => Delay1No503_out);

Delay1No504_out_to_Subtract32_5_impl_parent_implementedSystem_port_0_cast <= Delay1No504_out;
Delay1No505_out_to_Subtract32_5_impl_parent_implementedSystem_port_1_cast <= Delay1No505_out;
   Subtract32_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract32_5_impl_out,
                 X => Delay1No504_out_to_Subtract32_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No505_out_to_Subtract32_5_impl_parent_implementedSystem_port_1_cast);

SharedReg216_out_to_MUX_Subtract32_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg216_out;
SharedReg768_out_to_MUX_Subtract32_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg768_out;
SharedReg469_out_to_MUX_Subtract32_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg469_out;
SharedReg903_out_to_MUX_Subtract32_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg903_out;
SharedReg591_out_to_MUX_Subtract32_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg591_out;
SharedReg185_out_to_MUX_Subtract32_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg185_out;
SharedReg286_out_to_MUX_Subtract32_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg286_out;
SharedReg1029_out_to_MUX_Subtract32_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1029_out;
SharedReg662_out_to_MUX_Subtract32_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg662_out;
SharedReg317_out_to_MUX_Subtract32_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg317_out;
SharedReg13_out_to_MUX_Subtract32_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg13_out;
SharedReg12_out_to_MUX_Subtract32_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg12_out;
   MUX_Subtract32_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg216_out_to_MUX_Subtract32_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg768_out_to_MUX_Subtract32_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg13_out_to_MUX_Subtract32_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg12_out_to_MUX_Subtract32_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg469_out_to_MUX_Subtract32_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg903_out_to_MUX_Subtract32_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg591_out_to_MUX_Subtract32_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg185_out_to_MUX_Subtract32_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg286_out_to_MUX_Subtract32_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1029_out_to_MUX_Subtract32_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg662_out_to_MUX_Subtract32_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg317_out_to_MUX_Subtract32_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract32_5_impl_0_out);

   Delay1No504_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract32_5_impl_0_out,
                 Y => Delay1No504_out);

SharedReg315_out_to_MUX_Subtract32_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg315_out;
SharedReg466_out_to_MUX_Subtract32_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg466_out;
SharedReg998_out_to_MUX_Subtract32_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg998_out;
SharedReg975_out_to_MUX_Subtract32_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg975_out;
SharedReg464_out_to_MUX_Subtract32_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg464_out;
SharedReg150_out_to_MUX_Subtract32_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg150_out;
SharedReg289_out_to_MUX_Subtract32_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg289_out;
SharedReg1065_out_to_MUX_Subtract32_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1065_out;
SharedReg843_out_to_MUX_Subtract32_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg843_out;
SharedReg296_out_to_MUX_Subtract32_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg296_out;
SharedReg29_out_to_MUX_Subtract32_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg29_out;
SharedReg28_out_to_MUX_Subtract32_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg28_out;
   MUX_Subtract32_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg315_out_to_MUX_Subtract32_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg466_out_to_MUX_Subtract32_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg29_out_to_MUX_Subtract32_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg28_out_to_MUX_Subtract32_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg998_out_to_MUX_Subtract32_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg975_out_to_MUX_Subtract32_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg464_out_to_MUX_Subtract32_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg150_out_to_MUX_Subtract32_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg289_out_to_MUX_Subtract32_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1065_out_to_MUX_Subtract32_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg843_out_to_MUX_Subtract32_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg296_out_to_MUX_Subtract32_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract32_5_impl_1_out);

   Delay1No505_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract32_5_impl_1_out,
                 Y => Delay1No505_out);

Delay1No506_out_to_Subtract32_6_impl_parent_implementedSystem_port_0_cast <= Delay1No506_out;
Delay1No507_out_to_Subtract32_6_impl_parent_implementedSystem_port_1_cast <= Delay1No507_out;
   Subtract32_6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract32_6_impl_out,
                 X => Delay1No506_out_to_Subtract32_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No507_out_to_Subtract32_6_impl_parent_implementedSystem_port_1_cast);

SharedReg11_out_to_MUX_Subtract32_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg11_out;
SharedReg909_out_to_MUX_Subtract32_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg909_out;
SharedReg908_out_to_MUX_Subtract32_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg908_out;
SharedReg473_out_to_MUX_Subtract32_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg473_out;
SharedReg663_out_to_MUX_Subtract32_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg663_out;
SharedReg63_out_to_MUX_Subtract32_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg63_out;
SharedReg321_out_to_MUX_Subtract32_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg321_out;
SharedReg218_out_to_MUX_Subtract32_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg218_out;
SharedReg1034_out_to_MUX_Subtract32_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1034_out;
SharedReg665_out_to_MUX_Subtract32_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg665_out;
SharedReg703_out_to_MUX_Subtract32_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg703_out;
SharedReg6_out_to_MUX_Subtract32_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg6_out;
   MUX_Subtract32_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg11_out_to_MUX_Subtract32_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg909_out_to_MUX_Subtract32_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg703_out_to_MUX_Subtract32_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg6_out_to_MUX_Subtract32_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg908_out_to_MUX_Subtract32_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg473_out_to_MUX_Subtract32_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg663_out_to_MUX_Subtract32_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg63_out_to_MUX_Subtract32_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg321_out_to_MUX_Subtract32_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg218_out_to_MUX_Subtract32_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1034_out_to_MUX_Subtract32_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg665_out_to_MUX_Subtract32_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract32_6_impl_0_out);

   Delay1No506_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract32_6_impl_0_out,
                 Y => Delay1No506_out);

SharedReg27_out_to_MUX_Subtract32_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg27_out;
Delay5No48_out_to_MUX_Subtract32_6_impl_1_parent_implementedSystem_port_2_cast <= Delay5No48_out;
SharedReg979_out_to_MUX_Subtract32_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg979_out;
SharedReg872_out_to_MUX_Subtract32_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg872_out;
SharedReg845_out_to_MUX_Subtract32_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg845_out;
SharedReg355_out_to_MUX_Subtract32_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg355_out;
SharedReg389_out_to_MUX_Subtract32_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg389_out;
SharedReg222_out_to_MUX_Subtract32_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg222_out;
Delay12No20_out_to_MUX_Subtract32_6_impl_1_parent_implementedSystem_port_9_cast <= Delay12No20_out;
SharedReg847_out_to_MUX_Subtract32_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg847_out;
SharedReg479_out_to_MUX_Subtract32_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg479_out;
SharedReg22_out_to_MUX_Subtract32_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg22_out;
   MUX_Subtract32_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg27_out_to_MUX_Subtract32_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay5No48_out_to_MUX_Subtract32_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg479_out_to_MUX_Subtract32_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg22_out_to_MUX_Subtract32_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg979_out_to_MUX_Subtract32_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg872_out_to_MUX_Subtract32_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg845_out_to_MUX_Subtract32_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg355_out_to_MUX_Subtract32_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg389_out_to_MUX_Subtract32_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg222_out_to_MUX_Subtract32_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay12No20_out_to_MUX_Subtract32_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg847_out_to_MUX_Subtract32_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract32_6_impl_1_out);

   Delay1No507_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract32_6_impl_1_out,
                 Y => Delay1No507_out);

Delay1No508_out_to_Subtract43_0_impl_parent_implementedSystem_port_0_cast <= Delay1No508_out;
Delay1No509_out_to_Subtract43_0_impl_parent_implementedSystem_port_1_cast <= Delay1No509_out;
   Subtract43_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract43_0_impl_out,
                 X => Delay1No508_out_to_Subtract43_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No509_out_to_Subtract43_0_impl_parent_implementedSystem_port_1_cast);

SharedReg331_out_to_MUX_Subtract43_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg331_out;
SharedReg10_out_to_MUX_Subtract43_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg10_out;
SharedReg11_out_to_MUX_Subtract43_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg11_out;
SharedReg567_out_to_MUX_Subtract43_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg567_out;
SharedReg884_out_to_MUX_Subtract43_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg884_out;
SharedReg249_out_to_MUX_Subtract43_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg249_out;
SharedReg883_out_to_MUX_Subtract43_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg883_out;
SharedReg566_out_to_MUX_Subtract43_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg566_out;
SharedReg99_out_to_MUX_Subtract43_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg99_out;
SharedReg1004_out_to_MUX_Subtract43_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1004_out;
SharedReg1071_out_to_MUX_Subtract43_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1071_out;
SharedReg940_out_to_MUX_Subtract43_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg940_out;
   MUX_Subtract43_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg331_out_to_MUX_Subtract43_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg10_out_to_MUX_Subtract43_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1071_out_to_MUX_Subtract43_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg940_out_to_MUX_Subtract43_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg11_out_to_MUX_Subtract43_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg567_out_to_MUX_Subtract43_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg884_out_to_MUX_Subtract43_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg249_out_to_MUX_Subtract43_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg883_out_to_MUX_Subtract43_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg566_out_to_MUX_Subtract43_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg99_out_to_MUX_Subtract43_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1004_out_to_MUX_Subtract43_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract43_0_impl_0_out);

   Delay1No508_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract43_0_impl_0_out,
                 Y => Delay1No508_out);

SharedReg301_out_to_MUX_Subtract43_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg301_out;
SharedReg26_out_to_MUX_Subtract43_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg26_out;
SharedReg27_out_to_MUX_Subtract43_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg27_out;
SharedReg432_out_to_MUX_Subtract43_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg432_out;
SharedReg961_out_to_MUX_Subtract43_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg961_out;
SharedReg128_out_to_MUX_Subtract43_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg128_out;
SharedReg960_out_to_MUX_Subtract43_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg960_out;
SharedReg666_out_to_MUX_Subtract43_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg666_out;
SharedReg202_out_to_MUX_Subtract43_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg202_out;
SharedReg568_out_to_MUX_Subtract43_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg568_out;
SharedReg1074_out_to_MUX_Subtract43_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1074_out;
SharedReg960_out_to_MUX_Subtract43_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg960_out;
   MUX_Subtract43_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg301_out_to_MUX_Subtract43_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg26_out_to_MUX_Subtract43_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1074_out_to_MUX_Subtract43_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg960_out_to_MUX_Subtract43_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg27_out_to_MUX_Subtract43_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg432_out_to_MUX_Subtract43_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg961_out_to_MUX_Subtract43_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg128_out_to_MUX_Subtract43_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg960_out_to_MUX_Subtract43_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg666_out_to_MUX_Subtract43_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg202_out_to_MUX_Subtract43_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg568_out_to_MUX_Subtract43_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract43_0_impl_1_out);

   Delay1No509_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract43_0_impl_1_out,
                 Y => Delay1No509_out);

Delay1No510_out_to_Subtract44_6_impl_parent_implementedSystem_port_0_cast <= Delay1No510_out;
Delay1No511_out_to_Subtract44_6_impl_parent_implementedSystem_port_1_cast <= Delay1No511_out;
   Subtract44_6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract44_6_impl_out,
                 X => Delay1No510_out_to_Subtract44_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No511_out_to_Subtract44_6_impl_parent_implementedSystem_port_1_cast);

SharedReg12_out_to_MUX_Subtract44_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg12_out;
SharedReg600_out_to_MUX_Subtract44_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg600_out;
SharedReg477_out_to_MUX_Subtract44_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg477_out;
SharedReg218_out_to_MUX_Subtract44_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg218_out;
SharedReg907_out_to_MUX_Subtract44_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg907_out;
SharedReg598_out_to_MUX_Subtract44_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg598_out;
SharedReg702_out_to_MUX_Subtract44_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg702_out;
SharedReg1001_out_to_MUX_Subtract44_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1001_out;
SharedReg356_out_to_MUX_Subtract44_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg356_out;
SharedReg958_out_to_MUX_Subtract44_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg958_out;
SharedReg359_out_to_MUX_Subtract44_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg359_out;
SharedReg10_out_to_MUX_Subtract44_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg10_out;
   MUX_Subtract44_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg12_out_to_MUX_Subtract44_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg600_out_to_MUX_Subtract44_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg359_out_to_MUX_Subtract44_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg10_out_to_MUX_Subtract44_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg477_out_to_MUX_Subtract44_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg218_out_to_MUX_Subtract44_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg907_out_to_MUX_Subtract44_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg598_out_to_MUX_Subtract44_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg702_out_to_MUX_Subtract44_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1001_out_to_MUX_Subtract44_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg356_out_to_MUX_Subtract44_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg958_out_to_MUX_Subtract44_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract44_6_impl_0_out);

   Delay1No510_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract44_6_impl_0_out,
                 Y => Delay1No510_out);

SharedReg28_out_to_MUX_Subtract44_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg28_out;
SharedReg597_out_to_MUX_Subtract44_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg597_out;
SharedReg475_out_to_MUX_Subtract44_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg475_out;
SharedReg154_out_to_MUX_Subtract44_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg154_out;
SharedReg978_out_to_MUX_Subtract44_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg978_out;
SharedReg595_out_to_MUX_Subtract44_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg595_out;
SharedReg473_out_to_MUX_Subtract44_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg473_out;
SharedReg601_out_to_MUX_Subtract44_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg601_out;
SharedReg361_out_to_MUX_Subtract44_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg361_out;
SharedReg978_out_to_MUX_Subtract44_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg978_out;
SharedReg325_out_to_MUX_Subtract44_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg325_out;
SharedReg26_out_to_MUX_Subtract44_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg26_out;
   MUX_Subtract44_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg28_out_to_MUX_Subtract44_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg597_out_to_MUX_Subtract44_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg325_out_to_MUX_Subtract44_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg26_out_to_MUX_Subtract44_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg475_out_to_MUX_Subtract44_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg154_out_to_MUX_Subtract44_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg978_out_to_MUX_Subtract44_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg595_out_to_MUX_Subtract44_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg473_out_to_MUX_Subtract44_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg601_out_to_MUX_Subtract44_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg361_out_to_MUX_Subtract44_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg978_out_to_MUX_Subtract44_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract44_6_impl_1_out);

   Delay1No511_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract44_6_impl_1_out,
                 Y => Delay1No511_out);

Delay1No512_out_to_Subtract49_1_impl_parent_implementedSystem_port_0_cast <= Delay1No512_out;
Delay1No513_out_to_Subtract49_1_impl_parent_implementedSystem_port_1_cast <= Delay1No513_out;
   Subtract49_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract49_1_impl_out,
                 X => Delay1No512_out_to_Subtract49_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No513_out_to_Subtract49_1_impl_parent_implementedSystem_port_1_cast);

SharedReg165_out_to_MUX_Subtract49_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg165_out;
SharedReg943_out_to_MUX_Subtract49_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg943_out;
SharedReg375_out_to_MUX_Subtract49_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg375_out;
SharedReg10_out_to_MUX_Subtract49_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg10_out;
SharedReg11_out_to_MUX_Subtract49_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg11_out;
SharedReg104_out_to_MUX_Subtract49_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg104_out;
SharedReg780_out_to_MUX_Subtract49_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg780_out;
SharedReg573_out_to_MUX_Subtract49_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg573_out;
SharedReg339_out_to_MUX_Subtract49_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg339_out;
SharedReg72_out_to_MUX_Subtract49_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg72_out;
SharedReg441_out_to_MUX_Subtract49_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg441_out;
SharedReg335_out_to_MUX_Subtract49_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg335_out;
   MUX_Subtract49_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg165_out_to_MUX_Subtract49_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg943_out_to_MUX_Subtract49_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg441_out_to_MUX_Subtract49_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg335_out_to_MUX_Subtract49_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg375_out_to_MUX_Subtract49_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg10_out_to_MUX_Subtract49_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg11_out_to_MUX_Subtract49_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg104_out_to_MUX_Subtract49_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg780_out_to_MUX_Subtract49_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg573_out_to_MUX_Subtract49_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg339_out_to_MUX_Subtract49_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg72_out_to_MUX_Subtract49_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract49_1_impl_0_out);

   Delay1No512_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract49_1_impl_0_out,
                 Y => Delay1No512_out);

SharedReg378_out_to_MUX_Subtract49_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg378_out;
SharedReg963_out_to_MUX_Subtract49_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg963_out;
SharedReg259_out_to_MUX_Subtract49_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg259_out;
SharedReg26_out_to_MUX_Subtract49_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg26_out;
SharedReg27_out_to_MUX_Subtract49_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg27_out;
SharedReg256_out_to_MUX_Subtract49_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg256_out;
SharedReg777_out_to_MUX_Subtract49_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg777_out;
SharedReg985_out_to_MUX_Subtract49_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg985_out;
SharedReg236_out_to_MUX_Subtract49_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg236_out;
SharedReg41_out_to_MUX_Subtract49_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg41_out;
SharedReg984_out_to_MUX_Subtract49_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg984_out;
SharedReg258_out_to_MUX_Subtract49_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg258_out;
   MUX_Subtract49_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg378_out_to_MUX_Subtract49_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg963_out_to_MUX_Subtract49_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg984_out_to_MUX_Subtract49_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg258_out_to_MUX_Subtract49_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg259_out_to_MUX_Subtract49_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg26_out_to_MUX_Subtract49_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg27_out_to_MUX_Subtract49_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg256_out_to_MUX_Subtract49_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg777_out_to_MUX_Subtract49_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg985_out_to_MUX_Subtract49_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg236_out_to_MUX_Subtract49_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg41_out_to_MUX_Subtract49_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract49_1_impl_1_out);

   Delay1No513_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract49_1_impl_1_out,
                 Y => Delay1No513_out);

Delay1No514_out_to_Subtract116_6_impl_parent_implementedSystem_port_0_cast <= Delay1No514_out;
Delay1No515_out_to_Subtract116_6_impl_parent_implementedSystem_port_1_cast <= Delay1No515_out;
   Subtract116_6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract116_6_impl_out,
                 X => Delay1No514_out_to_Subtract116_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No515_out_to_Subtract116_6_impl_parent_implementedSystem_port_1_cast);

SharedReg14_out_to_MUX_Subtract116_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg14_out;
SharedReg157_out_to_MUX_Subtract116_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg157_out;
SharedReg874_out_to_MUX_Subtract116_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg874_out;
SharedReg703_out_to_MUX_Subtract116_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg703_out;
SharedReg360_out_to_MUX_Subtract116_6_impl_0_parent_implementedSystem_port_5_cast <= SharedReg360_out;
SharedReg94_out_to_MUX_Subtract116_6_impl_0_parent_implementedSystem_port_6_cast <= SharedReg94_out;
SharedReg126_out_to_MUX_Subtract116_6_impl_0_parent_implementedSystem_port_7_cast <= SharedReg126_out;
SharedReg320_out_to_MUX_Subtract116_6_impl_0_parent_implementedSystem_port_8_cast <= SharedReg320_out;
SharedReg1067_out_to_MUX_Subtract116_6_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1067_out;
SharedReg223_out_to_MUX_Subtract116_6_impl_0_parent_implementedSystem_port_10_cast <= SharedReg223_out;
SharedReg873_out_to_MUX_Subtract116_6_impl_0_parent_implementedSystem_port_11_cast <= SharedReg873_out;
SharedReg13_out_to_MUX_Subtract116_6_impl_0_parent_implementedSystem_port_12_cast <= SharedReg13_out;
   MUX_Subtract116_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg14_out_to_MUX_Subtract116_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg157_out_to_MUX_Subtract116_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg873_out_to_MUX_Subtract116_6_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg13_out_to_MUX_Subtract116_6_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg874_out_to_MUX_Subtract116_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg703_out_to_MUX_Subtract116_6_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg360_out_to_MUX_Subtract116_6_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg94_out_to_MUX_Subtract116_6_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg126_out_to_MUX_Subtract116_6_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg320_out_to_MUX_Subtract116_6_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1067_out_to_MUX_Subtract116_6_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg223_out_to_MUX_Subtract116_6_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract116_6_impl_0_out);

   Delay1No514_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract116_6_impl_0_out,
                 Y => Delay1No514_out);

SharedReg30_out_to_MUX_Subtract116_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg30_out;
SharedReg357_out_to_MUX_Subtract116_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg357_out;
SharedReg701_out_to_MUX_Subtract116_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg701_out;
SharedReg1002_out_to_MUX_Subtract116_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1002_out;
SharedReg189_out_to_MUX_Subtract116_6_impl_1_parent_implementedSystem_port_5_cast <= SharedReg189_out;
SharedReg381_out_to_MUX_Subtract116_6_impl_1_parent_implementedSystem_port_6_cast <= SharedReg381_out;
SharedReg187_out_to_MUX_Subtract116_6_impl_1_parent_implementedSystem_port_7_cast <= SharedReg187_out;
SharedReg324_out_to_MUX_Subtract116_6_impl_1_parent_implementedSystem_port_8_cast <= SharedReg324_out;
SharedReg1080_out_to_MUX_Subtract116_6_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1080_out;
SharedReg392_out_to_MUX_Subtract116_6_impl_1_parent_implementedSystem_port_10_cast <= SharedReg392_out;
SharedReg875_out_to_MUX_Subtract116_6_impl_1_parent_implementedSystem_port_11_cast <= SharedReg875_out;
SharedReg29_out_to_MUX_Subtract116_6_impl_1_parent_implementedSystem_port_12_cast <= SharedReg29_out;
   MUX_Subtract116_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg30_out_to_MUX_Subtract116_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg357_out_to_MUX_Subtract116_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg875_out_to_MUX_Subtract116_6_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg29_out_to_MUX_Subtract116_6_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg701_out_to_MUX_Subtract116_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1002_out_to_MUX_Subtract116_6_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg189_out_to_MUX_Subtract116_6_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg381_out_to_MUX_Subtract116_6_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg187_out_to_MUX_Subtract116_6_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg324_out_to_MUX_Subtract116_6_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1080_out_to_MUX_Subtract116_6_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg392_out_to_MUX_Subtract116_6_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract116_6_impl_1_out);

   Delay1No515_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract116_6_impl_1_out,
                 Y => Delay1No515_out);

Delay1No516_out_to_Subtract58_0_impl_parent_implementedSystem_port_0_cast <= Delay1No516_out;
Delay1No517_out_to_Subtract58_0_impl_parent_implementedSystem_port_1_cast <= Delay1No517_out;
   Subtract58_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract58_0_impl_out,
                 X => Delay1No516_out_to_Subtract58_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No517_out_to_Subtract58_0_impl_parent_implementedSystem_port_1_cast);

SharedReg852_out_to_MUX_Subtract58_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg852_out;
SharedReg13_out_to_MUX_Subtract58_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg13_out;
SharedReg12_out_to_MUX_Subtract58_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg12_out;
SharedReg129_out_to_MUX_Subtract58_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg129_out;
SharedReg435_out_to_MUX_Subtract58_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg435_out;
SharedReg669_out_to_MUX_Subtract58_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg669_out;
SharedReg332_out_to_MUX_Subtract58_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg332_out;
SharedReg68_out_to_MUX_Subtract58_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg68_out;
SharedReg433_out_to_MUX_Subtract58_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg433_out;
SharedReg326_out_to_MUX_Subtract58_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg326_out;
SharedReg159_out_to_MUX_Subtract58_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg159_out;
SharedReg253_out_to_MUX_Subtract58_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg253_out;
   MUX_Subtract58_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg852_out_to_MUX_Subtract58_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg13_out_to_MUX_Subtract58_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg159_out_to_MUX_Subtract58_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg253_out_to_MUX_Subtract58_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg12_out_to_MUX_Subtract58_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg129_out_to_MUX_Subtract58_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg435_out_to_MUX_Subtract58_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg669_out_to_MUX_Subtract58_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg332_out_to_MUX_Subtract58_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg68_out_to_MUX_Subtract58_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg433_out_to_MUX_Subtract58_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg326_out_to_MUX_Subtract58_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract58_0_impl_0_out);

   Delay1No516_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract58_0_impl_0_out,
                 Y => Delay1No516_out);

SharedReg671_out_to_MUX_Subtract58_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg671_out;
SharedReg29_out_to_MUX_Subtract58_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg29_out;
SharedReg28_out_to_MUX_Subtract58_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg28_out;
SharedReg298_out_to_MUX_Subtract58_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg298_out;
SharedReg432_out_to_MUX_Subtract58_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg432_out;
SharedReg982_out_to_MUX_Subtract58_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg982_out;
SharedReg203_out_to_MUX_Subtract58_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg203_out;
SharedReg158_out_to_MUX_Subtract58_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg158_out;
SharedReg1004_out_to_MUX_Subtract58_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1004_out;
SharedReg300_out_to_MUX_Subtract58_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg300_out;
SharedReg369_out_to_MUX_Subtract58_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg369_out;
SharedReg367_out_to_MUX_Subtract58_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg367_out;
   MUX_Subtract58_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg671_out_to_MUX_Subtract58_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg29_out_to_MUX_Subtract58_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg369_out_to_MUX_Subtract58_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg367_out_to_MUX_Subtract58_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg28_out_to_MUX_Subtract58_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg298_out_to_MUX_Subtract58_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg432_out_to_MUX_Subtract58_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg982_out_to_MUX_Subtract58_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg203_out_to_MUX_Subtract58_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg158_out_to_MUX_Subtract58_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1004_out_to_MUX_Subtract58_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg300_out_to_MUX_Subtract58_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount121_out,
                 oMux => MUX_Subtract58_0_impl_1_out);

   Delay1No517_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract58_0_impl_1_out,
                 Y => Delay1No517_out);

Delay1No518_out_to_Subtract125_6_impl_parent_implementedSystem_port_0_cast <= Delay1No518_out;
Delay1No519_out_to_Subtract125_6_impl_parent_implementedSystem_port_1_cast <= Delay1No519_out;
   Subtract125_6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract125_6_impl_out,
                 X => Delay1No518_out_to_Subtract125_6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No519_out_to_Subtract125_6_impl_parent_implementedSystem_port_1_cast);

SharedReg15_out_to_MUX_Subtract125_6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg15_out;
SharedReg476_out_to_MUX_Subtract125_6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg476_out;
SharedReg323_out_to_MUX_Subtract125_6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg323_out;
SharedReg382_out_to_MUX_Subtract125_6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg382_out;
   MUX_Subtract125_6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg15_out_to_MUX_Subtract125_6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg476_out_to_MUX_Subtract125_6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg323_out_to_MUX_Subtract125_6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg382_out_to_MUX_Subtract125_6_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => MUX_Subtract125_6_impl_0_LUT_out,
                 oMux => MUX_Subtract125_6_impl_0_out);

   Delay1No518_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract125_6_impl_0_out,
                 Y => Delay1No518_out);

SharedReg31_out_to_MUX_Subtract125_6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg31_out;
SharedReg383_out_to_MUX_Subtract125_6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg383_out;
SharedReg1033_out_to_MUX_Subtract125_6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1033_out;
SharedReg387_out_to_MUX_Subtract125_6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg387_out;
   MUX_Subtract125_6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg31_out_to_MUX_Subtract125_6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg383_out_to_MUX_Subtract125_6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1033_out_to_MUX_Subtract125_6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg387_out_to_MUX_Subtract125_6_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => MUX_Subtract125_6_impl_1_LUT_out,
                 oMux => MUX_Subtract125_6_impl_1_out);

   Delay1No519_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract125_6_impl_1_out,
                 Y => Delay1No519_out);
   Constant2_0_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant2_0_impl_out);
   Constant11_0_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant11_0_impl_out);
   Constant4_0_impl_instance: Constant_float_8_23_cosnpi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant4_0_impl_out);
   Constant13_0_impl_instance: Constant_float_8_23_sinnpi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant13_0_impl_out);
   Constant5_0_impl_instance: Constant_float_8_23_cosn3_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant5_0_impl_out);
   Constant14_0_impl_instance: Constant_float_8_23_sinn3_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant14_0_impl_out);
   Constant6_0_impl_instance: Constant_float_8_23_cosnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant6_0_impl_out);
   Constant15_0_impl_instance: Constant_float_8_23_sinnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant15_0_impl_out);
   Constant7_0_impl_instance: Constant_float_8_23_cosn5_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant7_0_impl_out);
   Constant16_0_impl_instance: Constant_float_8_23_sinn5_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant16_0_impl_out);
   Constant8_0_impl_instance: Constant_float_8_23_cosn3_mult_pi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant8_0_impl_out);
   Constant17_0_impl_instance: Constant_float_8_23_sinn3_mult_pi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant17_0_impl_out);
   Constant9_0_impl_instance: Constant_float_8_23_cosn7_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant9_0_impl_out);
   Constant18_0_impl_instance: Constant_float_8_23_sinn7_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant18_0_impl_out);
   Constant_0_impl_instance: Constant_float_8_23_cosnpi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant_0_impl_out);
   Constant1_0_impl_instance: Constant_float_8_23_sinnpi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant1_0_impl_out);

   Delay6No_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg504_out,
                 Y => Delay6No_out);

   Delay6No1_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg508_out,
                 Y => Delay6No1_out);

   Delay6No2_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg512_out,
                 Y => Delay6No2_out);

   Delay6No3_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg516_out,
                 Y => Delay6No3_out);

   Delay6No4_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg520_out,
                 Y => Delay6No4_out);

   Delay6No5_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg524_out,
                 Y => Delay6No5_out);

   Delay6No6_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg528_out,
                 Y => Delay6No6_out);

   Delay6No7_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg531_out,
                 Y => Delay6No7_out);

   Delay6No8_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg534_out,
                 Y => Delay6No8_out);

   Delay6No9_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg537_out,
                 Y => Delay6No9_out);

   Delay6No10_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg540_out,
                 Y => Delay6No10_out);

   Delay6No11_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg543_out,
                 Y => Delay6No11_out);

   Delay6No12_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg546_out,
                 Y => Delay6No12_out);

   Delay6No13_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg549_out,
                 Y => Delay6No13_out);

   Delay15No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg253_out,
                 Y => Delay15No_out);

   Delay15No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg238_out,
                 Y => Delay15No1_out);

   Delay15No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg243_out,
                 Y => Delay15No2_out);

   Delay15No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg144_out,
                 Y => Delay15No3_out);

   Delay15No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg149_out,
                 Y => Delay15No4_out);

   Delay15No5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg217_out,
                 Y => Delay15No5_out);

   Delay15No6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg223_out,
                 Y => Delay15No6_out);

   Delay10No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg174_out,
                 Y => Delay10No2_out);

   Delay10No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg181_out,
                 Y => Delay10No3_out);

   Delay4No168_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg647_out,
                 Y => Delay4No168_out);

   Delay4No169_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg650_out,
                 Y => Delay4No169_out);

   Delay4No170_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg653_out,
                 Y => Delay4No170_out);

   Delay4No171_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg656_out,
                 Y => Delay4No171_out);

   Delay4No172_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg659_out,
                 Y => Delay4No172_out);

   Delay4No173_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg662_out,
                 Y => Delay4No173_out);

   Delay4No174_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg665_out,
                 Y => Delay4No174_out);

   Delay4No182_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg802_out,
                 Y => Delay4No182_out);

   Delay4No183_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg805_out,
                 Y => Delay4No183_out);

   Delay4No184_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg808_out,
                 Y => Delay4No184_out);

   Delay4No185_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg811_out,
                 Y => Delay4No185_out);

   Delay4No186_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg814_out,
                 Y => Delay4No186_out);

   Delay4No187_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg817_out,
                 Y => Delay4No187_out);

   Delay4No188_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg820_out,
                 Y => Delay4No188_out);

   Delay4No210_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg397_out,
                 Y => Delay4No210_out);

   Delay4No211_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg400_out,
                 Y => Delay4No211_out);

   Delay4No212_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg403_out,
                 Y => Delay4No212_out);

   Delay4No213_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg406_out,
                 Y => Delay4No213_out);

   Delay4No214_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg409_out,
                 Y => Delay4No214_out);

   Delay4No215_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg412_out,
                 Y => Delay4No215_out);

   Delay4No216_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg415_out,
                 Y => Delay4No216_out);

   Delay4No217_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg417_out,
                 Y => Delay4No217_out);

   Delay4No218_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg419_out,
                 Y => Delay4No218_out);

   Delay4No219_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg421_out,
                 Y => Delay4No219_out);

   Delay4No220_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg423_out,
                 Y => Delay4No220_out);

   Delay4No221_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg425_out,
                 Y => Delay4No221_out);

   Delay4No222_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg427_out,
                 Y => Delay4No222_out);

   Delay4No223_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg429_out,
                 Y => Delay4No223_out);

   Delay4No224_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg482_out,
                 Y => Delay4No224_out);

   Delay4No225_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg485_out,
                 Y => Delay4No225_out);

   Delay4No226_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg488_out,
                 Y => Delay4No226_out);

   Delay4No227_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg491_out,
                 Y => Delay4No227_out);

   Delay4No228_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg494_out,
                 Y => Delay4No228_out);

   Delay4No229_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg497_out,
                 Y => Delay4No229_out);

   Delay4No230_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg500_out,
                 Y => Delay4No230_out);

   Delay3No238_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg551_out,
                 Y => Delay3No238_out);

   Delay3No239_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg553_out,
                 Y => Delay3No239_out);

   Delay3No240_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg555_out,
                 Y => Delay3No240_out);

   Delay3No241_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg557_out,
                 Y => Delay3No241_out);

   Delay3No242_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg559_out,
                 Y => Delay3No242_out);

   Delay3No243_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg561_out,
                 Y => Delay3No243_out);

   Delay3No244_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg563_out,
                 Y => Delay3No244_out);

   Delay4No259_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg941_out,
                 Y => Delay4No259_out);

   Delay4No260_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg944_out,
                 Y => Delay4No260_out);

   Delay4No261_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg947_out,
                 Y => Delay4No261_out);

   Delay4No262_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg950_out,
                 Y => Delay4No262_out);

   Delay4No263_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg953_out,
                 Y => Delay4No263_out);

   Delay4No264_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg956_out,
                 Y => Delay4No264_out);

   Delay4No265_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg959_out,
                 Y => Delay4No265_out);

   Delay4No266_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg962_out,
                 Y => Delay4No266_out);

   Delay4No267_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg965_out,
                 Y => Delay4No267_out);

   Delay4No268_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg968_out,
                 Y => Delay4No268_out);

   Delay4No269_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg971_out,
                 Y => Delay4No269_out);

   Delay4No270_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg974_out,
                 Y => Delay4No270_out);

   Delay4No271_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg977_out,
                 Y => Delay4No271_out);

   Delay4No272_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg980_out,
                 Y => Delay4No272_out);

   Delay12No14_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1041_out,
                 Y => Delay12No14_out);

   Delay12No15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1011_out,
                 Y => Delay12No15_out);

   Delay12No16_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg989_out,
                 Y => Delay12No16_out);

   Delay12No17_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg992_out,
                 Y => Delay12No17_out);

   Delay12No18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg996_out,
                 Y => Delay12No18_out);

   Delay12No19_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1032_out,
                 Y => Delay12No19_out);

   Delay12No20_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1069_out,
                 Y => Delay12No20_out);

   Delay6No42_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg824_out,
                 Y => Delay6No42_out);

   Delay6No43_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg828_out,
                 Y => Delay6No43_out);

   Delay6No44_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg832_out,
                 Y => Delay6No44_out);

   Delay6No45_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg836_out,
                 Y => Delay6No45_out);

   Delay6No46_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg840_out,
                 Y => Delay6No46_out);

   Delay6No47_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg844_out,
                 Y => Delay6No47_out);

   Delay6No48_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg848_out,
                 Y => Delay6No48_out);

   Delay5No42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg886_out,
                 Y => Delay5No42_out);

   Delay5No43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg890_out,
                 Y => Delay5No43_out);

   Delay5No44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg894_out,
                 Y => Delay5No44_out);

   Delay5No45_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg898_out,
                 Y => Delay5No45_out);

   Delay5No46_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg902_out,
                 Y => Delay5No46_out);

   Delay5No47_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg906_out,
                 Y => Delay5No47_out);

   Delay5No48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg910_out,
                 Y => Delay5No48_out);

   MUX_y0_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount121_out,
                 Output => MUX_y0_re_0_0_LUT_out);

   MUX_y0_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount121_out,
                 Output => MUX_y0_im_0_0_LUT_out);

   MUX_y1_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount121_out,
                 Output => MUX_y1_re_0_0_LUT_out);

   MUX_y1_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount121_out,
                 Output => MUX_y1_im_0_0_LUT_out);

   MUX_y2_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount121_out,
                 Output => MUX_y2_re_0_0_LUT_out);

   MUX_y2_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount121_out,
                 Output => MUX_y2_im_0_0_LUT_out);

   MUX_y3_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount121_out,
                 Output => MUX_y3_re_0_0_LUT_out);

   MUX_y3_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount121_out,
                 Output => MUX_y3_im_0_0_LUT_out);

   MUX_y4_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount121_out,
                 Output => MUX_y4_re_0_0_LUT_out);

   MUX_y4_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount121_out,
                 Output => MUX_y4_im_0_0_LUT_out);

   MUX_y5_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount121_out,
                 Output => MUX_y5_re_0_0_LUT_out);

   MUX_y5_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount121_out,
                 Output => MUX_y5_im_0_0_LUT_out);

   MUX_y6_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount121_out,
                 Output => MUX_y6_re_0_0_LUT_out);

   MUX_y6_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount121_out,
                 Output => MUX_y6_im_0_0_LUT_out);

   MUX_y7_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount121_out,
                 Output => MUX_y7_re_0_0_LUT_out);

   MUX_y7_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount121_out,
                 Output => MUX_y7_im_0_0_LUT_out);

   MUX_y8_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount121_out,
                 Output => MUX_y8_re_0_0_LUT_out);

   MUX_y8_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount121_out,
                 Output => MUX_y8_im_0_0_LUT_out);

   MUX_y9_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount121_out,
                 Output => MUX_y9_re_0_0_LUT_out);

   MUX_y9_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount121_out,
                 Output => MUX_y9_im_0_0_LUT_out);

   MUX_y10_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount121_out,
                 Output => MUX_y10_re_0_0_LUT_out);

   MUX_y10_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount121_out,
                 Output => MUX_y10_im_0_0_LUT_out);

   MUX_y11_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount121_out,
                 Output => MUX_y11_re_0_0_LUT_out);

   MUX_y11_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount121_out,
                 Output => MUX_y11_im_0_0_LUT_out);

   MUX_y12_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount121_out,
                 Output => MUX_y12_re_0_0_LUT_out);

   MUX_y12_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount121_out,
                 Output => MUX_y12_im_0_0_LUT_out);

   MUX_y13_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount121_out,
                 Output => MUX_y13_re_0_0_LUT_out);

   MUX_y13_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount121_out,
                 Output => MUX_y13_im_0_0_LUT_out);

   MUX_y14_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount121_out,
                 Output => MUX_y14_re_0_0_LUT_out);

   MUX_y14_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount121_out,
                 Output => MUX_y14_im_0_0_LUT_out);

   MUX_y15_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount121_out,
                 Output => MUX_y15_re_0_0_LUT_out);

   MUX_y15_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount121_out,
                 Output => MUX_y15_im_0_0_LUT_out);

   MUX_Add130_6_impl_0_LUT_instance: GenericLut_LUTData_MUX_Add130_6_impl_0_LUT_wIn_4_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount121_out,
                 Output => MUX_Add130_6_impl_0_LUT_out);

   MUX_Add130_6_impl_1_LUT_instance: GenericLut_LUTData_MUX_Add130_6_impl_1_LUT_wIn_4_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount121_out,
                 Output => MUX_Add130_6_impl_1_LUT_out);

   MUX_Subtract125_6_impl_0_LUT_instance: GenericLut_LUTData_MUX_Subtract125_6_impl_0_LUT_wIn_4_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount121_out,
                 Output => MUX_Subtract125_6_impl_0_LUT_out);

   MUX_Subtract125_6_impl_1_LUT_instance: GenericLut_LUTData_MUX_Subtract125_6_impl_1_LUT_wIn_4_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount121_out,
                 Output => MUX_Subtract125_6_impl_1_LUT_out);

   SharedReg_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x0_re_0_out,
                 Y => SharedReg_out);

   SharedReg1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x0_im_0_out,
                 Y => SharedReg1_out);

   SharedReg2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x1_re_0_out,
                 Y => SharedReg2_out);

   SharedReg3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x1_im_0_out,
                 Y => SharedReg3_out);

   SharedReg4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x2_re_0_out,
                 Y => SharedReg4_out);

   SharedReg5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x2_im_0_out,
                 Y => SharedReg5_out);

   SharedReg6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x3_re_0_out,
                 Y => SharedReg6_out);

   SharedReg7_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x3_im_0_out,
                 Y => SharedReg7_out);

   SharedReg8_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x4_re_0_out,
                 Y => SharedReg8_out);

   SharedReg9_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x4_im_0_out,
                 Y => SharedReg9_out);

   SharedReg10_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x5_re_0_out,
                 Y => SharedReg10_out);

   SharedReg11_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x5_im_0_out,
                 Y => SharedReg11_out);

   SharedReg12_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x6_re_0_out,
                 Y => SharedReg12_out);

   SharedReg13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x6_im_0_out,
                 Y => SharedReg13_out);

   SharedReg14_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x7_re_0_out,
                 Y => SharedReg14_out);

   SharedReg15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x7_im_0_out,
                 Y => SharedReg15_out);

   SharedReg16_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x8_re_0_out,
                 Y => SharedReg16_out);

   SharedReg17_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x8_im_0_out,
                 Y => SharedReg17_out);

   SharedReg18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x9_re_0_out,
                 Y => SharedReg18_out);

   SharedReg19_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x9_im_0_out,
                 Y => SharedReg19_out);

   SharedReg20_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x10_re_0_out,
                 Y => SharedReg20_out);

   SharedReg21_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x10_im_0_out,
                 Y => SharedReg21_out);

   SharedReg22_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x11_re_0_out,
                 Y => SharedReg22_out);

   SharedReg23_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x11_im_0_out,
                 Y => SharedReg23_out);

   SharedReg24_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x12_re_0_out,
                 Y => SharedReg24_out);

   SharedReg25_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x12_im_0_out,
                 Y => SharedReg25_out);

   SharedReg26_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x13_re_0_out,
                 Y => SharedReg26_out);

   SharedReg27_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x13_im_0_out,
                 Y => SharedReg27_out);

   SharedReg28_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x14_re_0_out,
                 Y => SharedReg28_out);

   SharedReg29_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x14_im_0_out,
                 Y => SharedReg29_out);

   SharedReg30_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x15_re_0_out,
                 Y => SharedReg30_out);

   SharedReg31_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x15_im_0_out,
                 Y => SharedReg31_out);

   SharedReg32_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_0_impl_out,
                 Y => SharedReg32_out);

   SharedReg33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg32_out,
                 Y => SharedReg33_out);

   SharedReg34_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg33_out,
                 Y => SharedReg34_out);

   SharedReg35_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg34_out,
                 Y => SharedReg35_out);

   SharedReg36_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg35_out,
                 Y => SharedReg36_out);

   SharedReg37_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg36_out,
                 Y => SharedReg37_out);

   SharedReg38_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_1_impl_out,
                 Y => SharedReg38_out);

   SharedReg39_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg38_out,
                 Y => SharedReg39_out);

   SharedReg40_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg39_out,
                 Y => SharedReg40_out);

   SharedReg41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_2_impl_out,
                 Y => SharedReg41_out);

   SharedReg42_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg41_out,
                 Y => SharedReg42_out);

   SharedReg43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg42_out,
                 Y => SharedReg43_out);

   SharedReg44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_3_impl_out,
                 Y => SharedReg44_out);

   SharedReg45_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg44_out,
                 Y => SharedReg45_out);

   SharedReg46_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg45_out,
                 Y => SharedReg46_out);

   SharedReg47_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg46_out,
                 Y => SharedReg47_out);

   SharedReg48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_4_impl_out,
                 Y => SharedReg48_out);

   SharedReg49_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg48_out,
                 Y => SharedReg49_out);

   SharedReg50_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg49_out,
                 Y => SharedReg50_out);

   SharedReg51_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg50_out,
                 Y => SharedReg51_out);

   SharedReg52_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_5_impl_out,
                 Y => SharedReg52_out);

   SharedReg53_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg52_out,
                 Y => SharedReg53_out);

   SharedReg54_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg53_out,
                 Y => SharedReg54_out);

   SharedReg55_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg54_out,
                 Y => SharedReg55_out);

   SharedReg56_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg55_out,
                 Y => SharedReg56_out);

   SharedReg57_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg56_out,
                 Y => SharedReg57_out);

   SharedReg58_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg57_out,
                 Y => SharedReg58_out);

   SharedReg59_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg58_out,
                 Y => SharedReg59_out);

   SharedReg60_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_6_impl_out,
                 Y => SharedReg60_out);

   SharedReg61_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg60_out,
                 Y => SharedReg61_out);

   SharedReg62_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg61_out,
                 Y => SharedReg62_out);

   SharedReg63_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg62_out,
                 Y => SharedReg63_out);

   SharedReg64_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg63_out,
                 Y => SharedReg64_out);

   SharedReg65_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_0_impl_out,
                 Y => SharedReg65_out);

   SharedReg66_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg65_out,
                 Y => SharedReg66_out);

   SharedReg67_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg66_out,
                 Y => SharedReg67_out);

   SharedReg68_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg67_out,
                 Y => SharedReg68_out);

   SharedReg69_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_1_impl_out,
                 Y => SharedReg69_out);

   SharedReg70_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg69_out,
                 Y => SharedReg70_out);

   SharedReg71_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg70_out,
                 Y => SharedReg71_out);

   SharedReg72_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg71_out,
                 Y => SharedReg72_out);

   SharedReg73_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_2_impl_out,
                 Y => SharedReg73_out);

   SharedReg74_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg73_out,
                 Y => SharedReg74_out);

   SharedReg75_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg74_out,
                 Y => SharedReg75_out);

   SharedReg76_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg75_out,
                 Y => SharedReg76_out);

   SharedReg77_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_3_impl_out,
                 Y => SharedReg77_out);

   SharedReg78_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg77_out,
                 Y => SharedReg78_out);

   SharedReg79_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg78_out,
                 Y => SharedReg79_out);

   SharedReg80_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg79_out,
                 Y => SharedReg80_out);

   SharedReg81_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_4_impl_out,
                 Y => SharedReg81_out);

   SharedReg82_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg81_out,
                 Y => SharedReg82_out);

   SharedReg83_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg82_out,
                 Y => SharedReg83_out);

   SharedReg84_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg83_out,
                 Y => SharedReg84_out);

   SharedReg85_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg84_out,
                 Y => SharedReg85_out);

   SharedReg86_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_5_impl_out,
                 Y => SharedReg86_out);

   SharedReg87_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg86_out,
                 Y => SharedReg87_out);

   SharedReg88_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg87_out,
                 Y => SharedReg88_out);

   SharedReg89_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg88_out,
                 Y => SharedReg89_out);

   SharedReg90_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg89_out,
                 Y => SharedReg90_out);

   SharedReg91_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_6_impl_out,
                 Y => SharedReg91_out);

   SharedReg92_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg91_out,
                 Y => SharedReg92_out);

   SharedReg93_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg92_out,
                 Y => SharedReg93_out);

   SharedReg94_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg93_out,
                 Y => SharedReg94_out);

   SharedReg95_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add3_0_impl_out,
                 Y => SharedReg95_out);

   SharedReg96_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg95_out,
                 Y => SharedReg96_out);

   SharedReg97_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg96_out,
                 Y => SharedReg97_out);

   SharedReg98_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg97_out,
                 Y => SharedReg98_out);

   SharedReg99_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg98_out,
                 Y => SharedReg99_out);

   SharedReg100_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add3_1_impl_out,
                 Y => SharedReg100_out);

   SharedReg101_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg100_out,
                 Y => SharedReg101_out);

   SharedReg102_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg101_out,
                 Y => SharedReg102_out);

   SharedReg103_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg102_out,
                 Y => SharedReg103_out);

   SharedReg104_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg103_out,
                 Y => SharedReg104_out);

   SharedReg105_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add3_2_impl_out,
                 Y => SharedReg105_out);

   SharedReg106_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg105_out,
                 Y => SharedReg106_out);

   SharedReg107_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg106_out,
                 Y => SharedReg107_out);

   SharedReg108_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg107_out,
                 Y => SharedReg108_out);

   SharedReg109_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg108_out,
                 Y => SharedReg109_out);

   SharedReg110_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add3_3_impl_out,
                 Y => SharedReg110_out);

   SharedReg111_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg110_out,
                 Y => SharedReg111_out);

   SharedReg112_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg111_out,
                 Y => SharedReg112_out);

   SharedReg113_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg112_out,
                 Y => SharedReg113_out);

   SharedReg114_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add3_4_impl_out,
                 Y => SharedReg114_out);

   SharedReg115_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg114_out,
                 Y => SharedReg115_out);

   SharedReg116_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg115_out,
                 Y => SharedReg116_out);

   SharedReg117_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg116_out,
                 Y => SharedReg117_out);

   SharedReg118_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add3_5_impl_out,
                 Y => SharedReg118_out);

   SharedReg119_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg118_out,
                 Y => SharedReg119_out);

   SharedReg120_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg119_out,
                 Y => SharedReg120_out);

   SharedReg121_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg120_out,
                 Y => SharedReg121_out);

   SharedReg122_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg121_out,
                 Y => SharedReg122_out);

   SharedReg123_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add3_6_impl_out,
                 Y => SharedReg123_out);

   SharedReg124_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg123_out,
                 Y => SharedReg124_out);

   SharedReg125_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg124_out,
                 Y => SharedReg125_out);

   SharedReg126_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg125_out,
                 Y => SharedReg126_out);

   SharedReg127_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add12_0_impl_out,
                 Y => SharedReg127_out);

   SharedReg128_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg127_out,
                 Y => SharedReg128_out);

   SharedReg129_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg128_out,
                 Y => SharedReg129_out);

   SharedReg130_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add12_1_impl_out,
                 Y => SharedReg130_out);

   SharedReg131_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg130_out,
                 Y => SharedReg131_out);

   SharedReg132_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg131_out,
                 Y => SharedReg132_out);

   SharedReg133_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg132_out,
                 Y => SharedReg133_out);

   SharedReg134_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add12_2_impl_out,
                 Y => SharedReg134_out);

   SharedReg135_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg134_out,
                 Y => SharedReg135_out);

   SharedReg136_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg135_out,
                 Y => SharedReg136_out);

   SharedReg137_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg136_out,
                 Y => SharedReg137_out);

   SharedReg138_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg137_out,
                 Y => SharedReg138_out);

   SharedReg139_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add12_3_impl_out,
                 Y => SharedReg139_out);

   SharedReg140_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg139_out,
                 Y => SharedReg140_out);

   SharedReg141_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg140_out,
                 Y => SharedReg141_out);

   SharedReg142_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg141_out,
                 Y => SharedReg142_out);

   SharedReg143_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg142_out,
                 Y => SharedReg143_out);

   SharedReg144_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg143_out,
                 Y => SharedReg144_out);

   SharedReg145_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add12_4_impl_out,
                 Y => SharedReg145_out);

   SharedReg146_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg145_out,
                 Y => SharedReg146_out);

   SharedReg147_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg146_out,
                 Y => SharedReg147_out);

   SharedReg148_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg147_out,
                 Y => SharedReg148_out);

   SharedReg149_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg148_out,
                 Y => SharedReg149_out);

   SharedReg150_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add12_5_impl_out,
                 Y => SharedReg150_out);

   SharedReg151_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg150_out,
                 Y => SharedReg151_out);

   SharedReg152_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg151_out,
                 Y => SharedReg152_out);

   SharedReg153_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add12_6_impl_out,
                 Y => SharedReg153_out);

   SharedReg154_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg153_out,
                 Y => SharedReg154_out);

   SharedReg155_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg154_out,
                 Y => SharedReg155_out);

   SharedReg156_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg155_out,
                 Y => SharedReg156_out);

   SharedReg157_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg156_out,
                 Y => SharedReg157_out);

   SharedReg158_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add5_1_impl_out,
                 Y => SharedReg158_out);

   SharedReg159_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg158_out,
                 Y => SharedReg159_out);

   SharedReg160_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg159_out,
                 Y => SharedReg160_out);

   SharedReg161_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg160_out,
                 Y => SharedReg161_out);

   SharedReg162_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg161_out,
                 Y => SharedReg162_out);

   SharedReg163_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg162_out,
                 Y => SharedReg163_out);

   SharedReg164_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add5_2_impl_out,
                 Y => SharedReg164_out);

   SharedReg165_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg164_out,
                 Y => SharedReg165_out);

   SharedReg166_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg165_out,
                 Y => SharedReg166_out);

   SharedReg167_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg166_out,
                 Y => SharedReg167_out);

   SharedReg168_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg167_out,
                 Y => SharedReg168_out);

   SharedReg169_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg168_out,
                 Y => SharedReg169_out);

   SharedReg170_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add5_3_impl_out,
                 Y => SharedReg170_out);

   SharedReg171_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg170_out,
                 Y => SharedReg171_out);

   SharedReg172_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg171_out,
                 Y => SharedReg172_out);

   SharedReg173_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg172_out,
                 Y => SharedReg173_out);

   SharedReg174_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg173_out,
                 Y => SharedReg174_out);

   SharedReg175_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add5_4_impl_out,
                 Y => SharedReg175_out);

   SharedReg176_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg175_out,
                 Y => SharedReg176_out);

   SharedReg177_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg176_out,
                 Y => SharedReg177_out);

   SharedReg178_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg177_out,
                 Y => SharedReg178_out);

   SharedReg179_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg178_out,
                 Y => SharedReg179_out);

   SharedReg180_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg179_out,
                 Y => SharedReg180_out);

   SharedReg181_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg180_out,
                 Y => SharedReg181_out);

   SharedReg182_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add14_5_impl_out,
                 Y => SharedReg182_out);

   SharedReg183_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg182_out,
                 Y => SharedReg183_out);

   SharedReg184_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg183_out,
                 Y => SharedReg184_out);

   SharedReg185_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg184_out,
                 Y => SharedReg185_out);

   SharedReg186_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg185_out,
                 Y => SharedReg186_out);

   SharedReg187_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add14_6_impl_out,
                 Y => SharedReg187_out);

   SharedReg188_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg187_out,
                 Y => SharedReg188_out);

   SharedReg189_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg188_out,
                 Y => SharedReg189_out);

   SharedReg190_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg189_out,
                 Y => SharedReg190_out);

   SharedReg191_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add6_4_impl_out,
                 Y => SharedReg191_out);

   SharedReg192_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg191_out,
                 Y => SharedReg192_out);

   SharedReg193_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg192_out,
                 Y => SharedReg193_out);

   SharedReg194_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg193_out,
                 Y => SharedReg194_out);

   SharedReg195_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg194_out,
                 Y => SharedReg195_out);

   SharedReg196_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg195_out,
                 Y => SharedReg196_out);

   SharedReg197_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg196_out,
                 Y => SharedReg197_out);

   SharedReg198_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add15_3_impl_out,
                 Y => SharedReg198_out);

   SharedReg199_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg198_out,
                 Y => SharedReg199_out);

   SharedReg200_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg199_out,
                 Y => SharedReg200_out);

   SharedReg201_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg200_out,
                 Y => SharedReg201_out);

   SharedReg202_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add8_0_impl_out,
                 Y => SharedReg202_out);

   SharedReg203_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg202_out,
                 Y => SharedReg203_out);

   SharedReg204_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg203_out,
                 Y => SharedReg204_out);

   SharedReg205_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg204_out,
                 Y => SharedReg205_out);

   SharedReg206_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add8_4_impl_out,
                 Y => SharedReg206_out);

   SharedReg207_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg206_out,
                 Y => SharedReg207_out);

   SharedReg208_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg207_out,
                 Y => SharedReg208_out);

   SharedReg209_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg208_out,
                 Y => SharedReg209_out);

   SharedReg210_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg209_out,
                 Y => SharedReg210_out);

   SharedReg211_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg210_out,
                 Y => SharedReg211_out);

   SharedReg212_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add8_5_impl_out,
                 Y => SharedReg212_out);

   SharedReg213_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg212_out,
                 Y => SharedReg213_out);

   SharedReg214_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg213_out,
                 Y => SharedReg214_out);

   SharedReg215_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg214_out,
                 Y => SharedReg215_out);

   SharedReg216_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg215_out,
                 Y => SharedReg216_out);

   SharedReg217_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg216_out,
                 Y => SharedReg217_out);

   SharedReg218_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add8_6_impl_out,
                 Y => SharedReg218_out);

   SharedReg219_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg218_out,
                 Y => SharedReg219_out);

   SharedReg220_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg219_out,
                 Y => SharedReg220_out);

   SharedReg221_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg220_out,
                 Y => SharedReg221_out);

   SharedReg222_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg221_out,
                 Y => SharedReg222_out);

   SharedReg223_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg222_out,
                 Y => SharedReg223_out);

   SharedReg224_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add10_6_impl_out,
                 Y => SharedReg224_out);

   SharedReg225_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg224_out,
                 Y => SharedReg225_out);

   SharedReg226_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg225_out,
                 Y => SharedReg226_out);

   SharedReg227_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg226_out,
                 Y => SharedReg227_out);

   SharedReg228_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg227_out,
                 Y => SharedReg228_out);

   SharedReg229_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg228_out,
                 Y => SharedReg229_out);

   SharedReg230_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg229_out,
                 Y => SharedReg230_out);

   SharedReg231_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg230_out,
                 Y => SharedReg231_out);

   SharedReg232_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg231_out,
                 Y => SharedReg232_out);

   SharedReg233_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg232_out,
                 Y => SharedReg233_out);

   SharedReg234_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add23_1_impl_out,
                 Y => SharedReg234_out);

   SharedReg235_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg234_out,
                 Y => SharedReg235_out);

   SharedReg236_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg235_out,
                 Y => SharedReg236_out);

   SharedReg237_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg236_out,
                 Y => SharedReg237_out);

   SharedReg238_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg237_out,
                 Y => SharedReg238_out);

   SharedReg239_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add23_2_impl_out,
                 Y => SharedReg239_out);

   SharedReg240_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg239_out,
                 Y => SharedReg240_out);

   SharedReg241_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg240_out,
                 Y => SharedReg241_out);

   SharedReg242_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg241_out,
                 Y => SharedReg242_out);

   SharedReg243_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg242_out,
                 Y => SharedReg243_out);

   SharedReg244_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add23_3_impl_out,
                 Y => SharedReg244_out);

   SharedReg245_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg244_out,
                 Y => SharedReg245_out);

   SharedReg246_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg245_out,
                 Y => SharedReg246_out);

   SharedReg247_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg246_out,
                 Y => SharedReg247_out);

   SharedReg248_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg247_out,
                 Y => SharedReg248_out);

   SharedReg249_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add113_0_impl_out,
                 Y => SharedReg249_out);

   SharedReg250_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg249_out,
                 Y => SharedReg250_out);

   SharedReg251_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg250_out,
                 Y => SharedReg251_out);

   SharedReg252_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg251_out,
                 Y => SharedReg252_out);

   SharedReg253_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg252_out,
                 Y => SharedReg253_out);

   SharedReg254_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add113_1_impl_out,
                 Y => SharedReg254_out);

   SharedReg255_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg254_out,
                 Y => SharedReg255_out);

   SharedReg256_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg255_out,
                 Y => SharedReg256_out);

   SharedReg257_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg256_out,
                 Y => SharedReg257_out);

   SharedReg258_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg257_out,
                 Y => SharedReg258_out);

   SharedReg259_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg258_out,
                 Y => SharedReg259_out);

   SharedReg260_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add113_2_impl_out,
                 Y => SharedReg260_out);

   SharedReg261_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg260_out,
                 Y => SharedReg261_out);

   SharedReg262_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg261_out,
                 Y => SharedReg262_out);

   SharedReg263_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg262_out,
                 Y => SharedReg263_out);

   SharedReg264_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg263_out,
                 Y => SharedReg264_out);

   SharedReg265_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg264_out,
                 Y => SharedReg265_out);

   SharedReg266_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add113_3_impl_out,
                 Y => SharedReg266_out);

   SharedReg267_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg266_out,
                 Y => SharedReg267_out);

   SharedReg268_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg267_out,
                 Y => SharedReg268_out);

   SharedReg269_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg268_out,
                 Y => SharedReg269_out);

   SharedReg270_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg269_out,
                 Y => SharedReg270_out);

   SharedReg271_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg270_out,
                 Y => SharedReg271_out);

   SharedReg272_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add113_4_impl_out,
                 Y => SharedReg272_out);

   SharedReg273_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg272_out,
                 Y => SharedReg273_out);

   SharedReg274_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg273_out,
                 Y => SharedReg274_out);

   SharedReg275_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg274_out,
                 Y => SharedReg275_out);

   SharedReg276_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg275_out,
                 Y => SharedReg276_out);

   SharedReg277_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg276_out,
                 Y => SharedReg277_out);

   SharedReg278_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add24_5_impl_out,
                 Y => SharedReg278_out);

   SharedReg279_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg278_out,
                 Y => SharedReg279_out);

   SharedReg280_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg279_out,
                 Y => SharedReg280_out);

   SharedReg281_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg280_out,
                 Y => SharedReg281_out);

   SharedReg282_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg281_out,
                 Y => SharedReg282_out);

   SharedReg283_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg282_out,
                 Y => SharedReg283_out);

   SharedReg284_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg283_out,
                 Y => SharedReg284_out);

   SharedReg285_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg284_out,
                 Y => SharedReg285_out);

   SharedReg286_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add32_5_impl_out,
                 Y => SharedReg286_out);

   SharedReg287_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg286_out,
                 Y => SharedReg287_out);

   SharedReg288_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg287_out,
                 Y => SharedReg288_out);

   SharedReg289_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg288_out,
                 Y => SharedReg289_out);

   SharedReg290_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add122_5_impl_out,
                 Y => SharedReg290_out);

   SharedReg291_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg290_out,
                 Y => SharedReg291_out);

   SharedReg292_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg291_out,
                 Y => SharedReg292_out);

   SharedReg293_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg292_out,
                 Y => SharedReg293_out);

   SharedReg294_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg293_out,
                 Y => SharedReg294_out);

   SharedReg295_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg294_out,
                 Y => SharedReg295_out);

   SharedReg296_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg295_out,
                 Y => SharedReg296_out);

   SharedReg297_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add33_0_impl_out,
                 Y => SharedReg297_out);

   SharedReg298_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg297_out,
                 Y => SharedReg298_out);

   SharedReg299_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg298_out,
                 Y => SharedReg299_out);

   SharedReg300_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg299_out,
                 Y => SharedReg300_out);

   SharedReg301_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg300_out,
                 Y => SharedReg301_out);

   SharedReg302_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add33_2_impl_out,
                 Y => SharedReg302_out);

   SharedReg303_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg302_out,
                 Y => SharedReg303_out);

   SharedReg304_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg303_out,
                 Y => SharedReg304_out);

   SharedReg305_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg304_out,
                 Y => SharedReg305_out);

   SharedReg306_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg305_out,
                 Y => SharedReg306_out);

   SharedReg307_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg306_out,
                 Y => SharedReg307_out);

   SharedReg308_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add33_4_impl_out,
                 Y => SharedReg308_out);

   SharedReg309_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg308_out,
                 Y => SharedReg309_out);

   SharedReg310_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg309_out,
                 Y => SharedReg310_out);

   SharedReg311_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg310_out,
                 Y => SharedReg311_out);

   SharedReg312_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg311_out,
                 Y => SharedReg312_out);

   SharedReg313_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add33_5_impl_out,
                 Y => SharedReg313_out);

   SharedReg314_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg313_out,
                 Y => SharedReg314_out);

   SharedReg315_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg314_out,
                 Y => SharedReg315_out);

   SharedReg316_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg315_out,
                 Y => SharedReg316_out);

   SharedReg317_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg316_out,
                 Y => SharedReg317_out);

   SharedReg318_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg317_out,
                 Y => SharedReg318_out);

   SharedReg319_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg318_out,
                 Y => SharedReg319_out);

   SharedReg320_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add33_6_impl_out,
                 Y => SharedReg320_out);

   SharedReg321_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg320_out,
                 Y => SharedReg321_out);

   SharedReg322_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg321_out,
                 Y => SharedReg322_out);

   SharedReg323_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg322_out,
                 Y => SharedReg323_out);

   SharedReg324_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg323_out,
                 Y => SharedReg324_out);

   SharedReg325_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg324_out,
                 Y => SharedReg325_out);

   SharedReg326_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add123_0_impl_out,
                 Y => SharedReg326_out);

   SharedReg327_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg326_out,
                 Y => SharedReg327_out);

   SharedReg328_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg327_out,
                 Y => SharedReg328_out);

   SharedReg329_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg328_out,
                 Y => SharedReg329_out);

   SharedReg330_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg329_out,
                 Y => SharedReg330_out);

   SharedReg331_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg330_out,
                 Y => SharedReg331_out);

   SharedReg332_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg331_out,
                 Y => SharedReg332_out);

   SharedReg333_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg332_out,
                 Y => SharedReg333_out);

   SharedReg334_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg333_out,
                 Y => SharedReg334_out);

   SharedReg335_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add123_1_impl_out,
                 Y => SharedReg335_out);

   SharedReg336_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg335_out,
                 Y => SharedReg336_out);

   SharedReg337_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg336_out,
                 Y => SharedReg337_out);

   SharedReg338_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg337_out,
                 Y => SharedReg338_out);

   SharedReg339_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg338_out,
                 Y => SharedReg339_out);

   SharedReg340_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg339_out,
                 Y => SharedReg340_out);

   SharedReg341_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg340_out,
                 Y => SharedReg341_out);

   SharedReg342_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add123_2_impl_out,
                 Y => SharedReg342_out);

   SharedReg343_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg342_out,
                 Y => SharedReg343_out);

   SharedReg344_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg343_out,
                 Y => SharedReg344_out);

   SharedReg345_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg344_out,
                 Y => SharedReg345_out);

   SharedReg346_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg345_out,
                 Y => SharedReg346_out);

   SharedReg347_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg346_out,
                 Y => SharedReg347_out);

   SharedReg348_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg347_out,
                 Y => SharedReg348_out);

   SharedReg349_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg348_out,
                 Y => SharedReg349_out);

   SharedReg350_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add123_3_impl_out,
                 Y => SharedReg350_out);

   SharedReg351_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg350_out,
                 Y => SharedReg351_out);

   SharedReg352_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg351_out,
                 Y => SharedReg352_out);

   SharedReg353_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg352_out,
                 Y => SharedReg353_out);

   SharedReg354_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg353_out,
                 Y => SharedReg354_out);

   SharedReg355_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add123_6_impl_out,
                 Y => SharedReg355_out);

   SharedReg356_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg355_out,
                 Y => SharedReg356_out);

   SharedReg357_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg356_out,
                 Y => SharedReg357_out);

   SharedReg358_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg357_out,
                 Y => SharedReg358_out);

   SharedReg359_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg358_out,
                 Y => SharedReg359_out);

   SharedReg360_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg359_out,
                 Y => SharedReg360_out);

   SharedReg361_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg360_out,
                 Y => SharedReg361_out);

   SharedReg362_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg361_out,
                 Y => SharedReg362_out);

   SharedReg363_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add35_0_impl_out,
                 Y => SharedReg363_out);

   SharedReg364_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg363_out,
                 Y => SharedReg364_out);

   SharedReg365_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg364_out,
                 Y => SharedReg365_out);

   SharedReg366_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg365_out,
                 Y => SharedReg366_out);

   SharedReg367_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg366_out,
                 Y => SharedReg367_out);

   SharedReg368_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg367_out,
                 Y => SharedReg368_out);

   SharedReg369_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg368_out,
                 Y => SharedReg369_out);

   SharedReg370_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg369_out,
                 Y => SharedReg370_out);

   SharedReg371_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg370_out,
                 Y => SharedReg371_out);

   SharedReg372_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add35_1_impl_out,
                 Y => SharedReg372_out);

   SharedReg373_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg372_out,
                 Y => SharedReg373_out);

   SharedReg374_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg373_out,
                 Y => SharedReg374_out);

   SharedReg375_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg374_out,
                 Y => SharedReg375_out);

   SharedReg376_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg375_out,
                 Y => SharedReg376_out);

   SharedReg377_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg376_out,
                 Y => SharedReg377_out);

   SharedReg378_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg377_out,
                 Y => SharedReg378_out);

   SharedReg379_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg378_out,
                 Y => SharedReg379_out);

   SharedReg380_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg379_out,
                 Y => SharedReg380_out);

   SharedReg381_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add35_6_impl_out,
                 Y => SharedReg381_out);

   SharedReg382_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg381_out,
                 Y => SharedReg382_out);

   SharedReg383_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg382_out,
                 Y => SharedReg383_out);

   SharedReg384_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg383_out,
                 Y => SharedReg384_out);

   SharedReg385_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg384_out,
                 Y => SharedReg385_out);

   SharedReg386_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg385_out,
                 Y => SharedReg386_out);

   SharedReg387_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg386_out,
                 Y => SharedReg387_out);

   SharedReg388_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg387_out,
                 Y => SharedReg388_out);

   SharedReg389_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add130_6_impl_out,
                 Y => SharedReg389_out);

   SharedReg390_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg389_out,
                 Y => SharedReg390_out);

   SharedReg391_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg390_out,
                 Y => SharedReg391_out);

   SharedReg392_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg391_out,
                 Y => SharedReg392_out);

   SharedReg393_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg392_out,
                 Y => SharedReg393_out);

   SharedReg394_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg393_out,
                 Y => SharedReg394_out);

   SharedReg395_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_0_impl_out,
                 Y => SharedReg395_out);

   SharedReg396_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg395_out,
                 Y => SharedReg396_out);

   SharedReg397_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg396_out,
                 Y => SharedReg397_out);

   SharedReg398_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_1_impl_out,
                 Y => SharedReg398_out);

   SharedReg399_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg398_out,
                 Y => SharedReg399_out);

   SharedReg400_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg399_out,
                 Y => SharedReg400_out);

   SharedReg401_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_2_impl_out,
                 Y => SharedReg401_out);

   SharedReg402_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg401_out,
                 Y => SharedReg402_out);

   SharedReg403_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg402_out,
                 Y => SharedReg403_out);

   SharedReg404_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_3_impl_out,
                 Y => SharedReg404_out);

   SharedReg405_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg404_out,
                 Y => SharedReg405_out);

   SharedReg406_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg405_out,
                 Y => SharedReg406_out);

   SharedReg407_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_4_impl_out,
                 Y => SharedReg407_out);

   SharedReg408_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg407_out,
                 Y => SharedReg408_out);

   SharedReg409_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg408_out,
                 Y => SharedReg409_out);

   SharedReg410_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_5_impl_out,
                 Y => SharedReg410_out);

   SharedReg411_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg410_out,
                 Y => SharedReg411_out);

   SharedReg412_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg411_out,
                 Y => SharedReg412_out);

   SharedReg413_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_6_impl_out,
                 Y => SharedReg413_out);

   SharedReg414_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg413_out,
                 Y => SharedReg414_out);

   SharedReg415_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg414_out,
                 Y => SharedReg415_out);

   SharedReg416_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_0_impl_out,
                 Y => SharedReg416_out);

   SharedReg417_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg416_out,
                 Y => SharedReg417_out);

   SharedReg418_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_1_impl_out,
                 Y => SharedReg418_out);

   SharedReg419_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg418_out,
                 Y => SharedReg419_out);

   SharedReg420_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_2_impl_out,
                 Y => SharedReg420_out);

   SharedReg421_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg420_out,
                 Y => SharedReg421_out);

   SharedReg422_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_3_impl_out,
                 Y => SharedReg422_out);

   SharedReg423_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg422_out,
                 Y => SharedReg423_out);

   SharedReg424_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_4_impl_out,
                 Y => SharedReg424_out);

   SharedReg425_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg424_out,
                 Y => SharedReg425_out);

   SharedReg426_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_5_impl_out,
                 Y => SharedReg426_out);

   SharedReg427_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg426_out,
                 Y => SharedReg427_out);

   SharedReg428_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_6_impl_out,
                 Y => SharedReg428_out);

   SharedReg429_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg428_out,
                 Y => SharedReg429_out);

   SharedReg430_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_0_impl_out,
                 Y => SharedReg430_out);

   SharedReg431_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg430_out,
                 Y => SharedReg431_out);

   SharedReg432_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg431_out,
                 Y => SharedReg432_out);

   SharedReg433_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg432_out,
                 Y => SharedReg433_out);

   SharedReg434_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg433_out,
                 Y => SharedReg434_out);

   SharedReg435_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg434_out,
                 Y => SharedReg435_out);

   SharedReg436_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg435_out,
                 Y => SharedReg436_out);

   SharedReg437_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg436_out,
                 Y => SharedReg437_out);

   SharedReg438_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_1_impl_out,
                 Y => SharedReg438_out);

   SharedReg439_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg438_out,
                 Y => SharedReg439_out);

   SharedReg440_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg439_out,
                 Y => SharedReg440_out);

   SharedReg441_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg440_out,
                 Y => SharedReg441_out);

   SharedReg442_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg441_out,
                 Y => SharedReg442_out);

   SharedReg443_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg442_out,
                 Y => SharedReg443_out);

   SharedReg444_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg443_out,
                 Y => SharedReg444_out);

   SharedReg445_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_2_impl_out,
                 Y => SharedReg445_out);

   SharedReg446_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg445_out,
                 Y => SharedReg446_out);

   SharedReg447_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg446_out,
                 Y => SharedReg447_out);

   SharedReg448_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg447_out,
                 Y => SharedReg448_out);

   SharedReg449_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg448_out,
                 Y => SharedReg449_out);

   SharedReg450_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg449_out,
                 Y => SharedReg450_out);

   SharedReg451_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_3_impl_out,
                 Y => SharedReg451_out);

   SharedReg452_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg451_out,
                 Y => SharedReg452_out);

   SharedReg453_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg452_out,
                 Y => SharedReg453_out);

   SharedReg454_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg453_out,
                 Y => SharedReg454_out);

   SharedReg455_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg454_out,
                 Y => SharedReg455_out);

   SharedReg456_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg455_out,
                 Y => SharedReg456_out);

   SharedReg457_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg456_out,
                 Y => SharedReg457_out);

   SharedReg458_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_4_impl_out,
                 Y => SharedReg458_out);

   SharedReg459_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg458_out,
                 Y => SharedReg459_out);

   SharedReg460_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg459_out,
                 Y => SharedReg460_out);

   SharedReg461_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg460_out,
                 Y => SharedReg461_out);

   SharedReg462_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg461_out,
                 Y => SharedReg462_out);

   SharedReg463_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg462_out,
                 Y => SharedReg463_out);

   SharedReg464_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_5_impl_out,
                 Y => SharedReg464_out);

   SharedReg465_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg464_out,
                 Y => SharedReg465_out);

   SharedReg466_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg465_out,
                 Y => SharedReg466_out);

   SharedReg467_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg466_out,
                 Y => SharedReg467_out);

   SharedReg468_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg467_out,
                 Y => SharedReg468_out);

   SharedReg469_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg468_out,
                 Y => SharedReg469_out);

   SharedReg470_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg469_out,
                 Y => SharedReg470_out);

   SharedReg471_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg470_out,
                 Y => SharedReg471_out);

   SharedReg472_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg471_out,
                 Y => SharedReg472_out);

   SharedReg473_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_6_impl_out,
                 Y => SharedReg473_out);

   SharedReg474_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg473_out,
                 Y => SharedReg474_out);

   SharedReg475_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg474_out,
                 Y => SharedReg475_out);

   SharedReg476_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg475_out,
                 Y => SharedReg476_out);

   SharedReg477_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg476_out,
                 Y => SharedReg477_out);

   SharedReg478_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg477_out,
                 Y => SharedReg478_out);

   SharedReg479_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg478_out,
                 Y => SharedReg479_out);

   SharedReg480_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product5_0_impl_out,
                 Y => SharedReg480_out);

   SharedReg481_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg480_out,
                 Y => SharedReg481_out);

   SharedReg482_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg481_out,
                 Y => SharedReg482_out);

   SharedReg483_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product5_1_impl_out,
                 Y => SharedReg483_out);

   SharedReg484_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg483_out,
                 Y => SharedReg484_out);

   SharedReg485_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg484_out,
                 Y => SharedReg485_out);

   SharedReg486_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product5_2_impl_out,
                 Y => SharedReg486_out);

   SharedReg487_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg486_out,
                 Y => SharedReg487_out);

   SharedReg488_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg487_out,
                 Y => SharedReg488_out);

   SharedReg489_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product5_3_impl_out,
                 Y => SharedReg489_out);

   SharedReg490_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg489_out,
                 Y => SharedReg490_out);

   SharedReg491_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg490_out,
                 Y => SharedReg491_out);

   SharedReg492_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product5_4_impl_out,
                 Y => SharedReg492_out);

   SharedReg493_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg492_out,
                 Y => SharedReg493_out);

   SharedReg494_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg493_out,
                 Y => SharedReg494_out);

   SharedReg495_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product5_5_impl_out,
                 Y => SharedReg495_out);

   SharedReg496_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg495_out,
                 Y => SharedReg496_out);

   SharedReg497_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg496_out,
                 Y => SharedReg497_out);

   SharedReg498_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product5_6_impl_out,
                 Y => SharedReg498_out);

   SharedReg499_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg498_out,
                 Y => SharedReg499_out);

   SharedReg500_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg499_out,
                 Y => SharedReg500_out);

   SharedReg501_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product12_0_impl_out,
                 Y => SharedReg501_out);

   SharedReg502_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg501_out,
                 Y => SharedReg502_out);

   SharedReg503_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg502_out,
                 Y => SharedReg503_out);

   SharedReg504_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg503_out,
                 Y => SharedReg504_out);

   SharedReg505_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product12_1_impl_out,
                 Y => SharedReg505_out);

   SharedReg506_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg505_out,
                 Y => SharedReg506_out);

   SharedReg507_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg506_out,
                 Y => SharedReg507_out);

   SharedReg508_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg507_out,
                 Y => SharedReg508_out);

   SharedReg509_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product12_2_impl_out,
                 Y => SharedReg509_out);

   SharedReg510_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg509_out,
                 Y => SharedReg510_out);

   SharedReg511_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg510_out,
                 Y => SharedReg511_out);

   SharedReg512_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg511_out,
                 Y => SharedReg512_out);

   SharedReg513_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product12_3_impl_out,
                 Y => SharedReg513_out);

   SharedReg514_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg513_out,
                 Y => SharedReg514_out);

   SharedReg515_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg514_out,
                 Y => SharedReg515_out);

   SharedReg516_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg515_out,
                 Y => SharedReg516_out);

   SharedReg517_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product12_4_impl_out,
                 Y => SharedReg517_out);

   SharedReg518_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg517_out,
                 Y => SharedReg518_out);

   SharedReg519_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg518_out,
                 Y => SharedReg519_out);

   SharedReg520_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg519_out,
                 Y => SharedReg520_out);

   SharedReg521_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product12_5_impl_out,
                 Y => SharedReg521_out);

   SharedReg522_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg521_out,
                 Y => SharedReg522_out);

   SharedReg523_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg522_out,
                 Y => SharedReg523_out);

   SharedReg524_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg523_out,
                 Y => SharedReg524_out);

   SharedReg525_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product12_6_impl_out,
                 Y => SharedReg525_out);

   SharedReg526_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg525_out,
                 Y => SharedReg526_out);

   SharedReg527_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg526_out,
                 Y => SharedReg527_out);

   SharedReg528_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg527_out,
                 Y => SharedReg528_out);

   SharedReg529_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product22_0_impl_out,
                 Y => SharedReg529_out);

   SharedReg530_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg529_out,
                 Y => SharedReg530_out);

   SharedReg531_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg530_out,
                 Y => SharedReg531_out);

   SharedReg532_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product22_1_impl_out,
                 Y => SharedReg532_out);

   SharedReg533_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg532_out,
                 Y => SharedReg533_out);

   SharedReg534_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg533_out,
                 Y => SharedReg534_out);

   SharedReg535_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product22_2_impl_out,
                 Y => SharedReg535_out);

   SharedReg536_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg535_out,
                 Y => SharedReg536_out);

   SharedReg537_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg536_out,
                 Y => SharedReg537_out);

   SharedReg538_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product22_3_impl_out,
                 Y => SharedReg538_out);

   SharedReg539_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg538_out,
                 Y => SharedReg539_out);

   SharedReg540_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg539_out,
                 Y => SharedReg540_out);

   SharedReg541_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product22_4_impl_out,
                 Y => SharedReg541_out);

   SharedReg542_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg541_out,
                 Y => SharedReg542_out);

   SharedReg543_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg542_out,
                 Y => SharedReg543_out);

   SharedReg544_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product22_5_impl_out,
                 Y => SharedReg544_out);

   SharedReg545_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg544_out,
                 Y => SharedReg545_out);

   SharedReg546_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg545_out,
                 Y => SharedReg546_out);

   SharedReg547_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product22_6_impl_out,
                 Y => SharedReg547_out);

   SharedReg548_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg547_out,
                 Y => SharedReg548_out);

   SharedReg549_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg548_out,
                 Y => SharedReg549_out);

   SharedReg550_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_0_impl_out,
                 Y => SharedReg550_out);

   SharedReg551_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg550_out,
                 Y => SharedReg551_out);

   SharedReg552_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_1_impl_out,
                 Y => SharedReg552_out);

   SharedReg553_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg552_out,
                 Y => SharedReg553_out);

   SharedReg554_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_2_impl_out,
                 Y => SharedReg554_out);

   SharedReg555_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg554_out,
                 Y => SharedReg555_out);

   SharedReg556_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_3_impl_out,
                 Y => SharedReg556_out);

   SharedReg557_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg556_out,
                 Y => SharedReg557_out);

   SharedReg558_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_4_impl_out,
                 Y => SharedReg558_out);

   SharedReg559_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg558_out,
                 Y => SharedReg559_out);

   SharedReg560_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_5_impl_out,
                 Y => SharedReg560_out);

   SharedReg561_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg560_out,
                 Y => SharedReg561_out);

   SharedReg562_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_6_impl_out,
                 Y => SharedReg562_out);

   SharedReg563_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg562_out,
                 Y => SharedReg563_out);

   SharedReg564_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract3_0_impl_out,
                 Y => SharedReg564_out);

   SharedReg565_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg564_out,
                 Y => SharedReg565_out);

   SharedReg566_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg565_out,
                 Y => SharedReg566_out);

   SharedReg567_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg566_out,
                 Y => SharedReg567_out);

   SharedReg568_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg567_out,
                 Y => SharedReg568_out);

   SharedReg569_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg568_out,
                 Y => SharedReg569_out);

   SharedReg570_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract3_1_impl_out,
                 Y => SharedReg570_out);

   SharedReg571_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg570_out,
                 Y => SharedReg571_out);

   SharedReg572_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg571_out,
                 Y => SharedReg572_out);

   SharedReg573_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg572_out,
                 Y => SharedReg573_out);

   SharedReg574_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg573_out,
                 Y => SharedReg574_out);

   SharedReg575_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg574_out,
                 Y => SharedReg575_out);

   SharedReg576_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract3_2_impl_out,
                 Y => SharedReg576_out);

   SharedReg577_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg576_out,
                 Y => SharedReg577_out);

   SharedReg578_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg577_out,
                 Y => SharedReg578_out);

   SharedReg579_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg578_out,
                 Y => SharedReg579_out);

   SharedReg580_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract3_3_impl_out,
                 Y => SharedReg580_out);

   SharedReg581_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg580_out,
                 Y => SharedReg581_out);

   SharedReg582_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg581_out,
                 Y => SharedReg582_out);

   SharedReg583_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg582_out,
                 Y => SharedReg583_out);

   SharedReg584_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract3_4_impl_out,
                 Y => SharedReg584_out);

   SharedReg585_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg584_out,
                 Y => SharedReg585_out);

   SharedReg586_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg585_out,
                 Y => SharedReg586_out);

   SharedReg587_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg586_out,
                 Y => SharedReg587_out);

   SharedReg588_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg587_out,
                 Y => SharedReg588_out);

   SharedReg589_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract3_5_impl_out,
                 Y => SharedReg589_out);

   SharedReg590_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg589_out,
                 Y => SharedReg590_out);

   SharedReg591_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg590_out,
                 Y => SharedReg591_out);

   SharedReg592_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg591_out,
                 Y => SharedReg592_out);

   SharedReg593_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg592_out,
                 Y => SharedReg593_out);

   SharedReg594_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg593_out,
                 Y => SharedReg594_out);

   SharedReg595_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract3_6_impl_out,
                 Y => SharedReg595_out);

   SharedReg596_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg595_out,
                 Y => SharedReg596_out);

   SharedReg597_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg596_out,
                 Y => SharedReg597_out);

   SharedReg598_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg597_out,
                 Y => SharedReg598_out);

   SharedReg599_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg598_out,
                 Y => SharedReg599_out);

   SharedReg600_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg599_out,
                 Y => SharedReg600_out);

   SharedReg601_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg600_out,
                 Y => SharedReg601_out);

   SharedReg602_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg601_out,
                 Y => SharedReg602_out);

   SharedReg603_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product6_0_impl_out,
                 Y => SharedReg603_out);

   SharedReg604_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg603_out,
                 Y => SharedReg604_out);

   SharedReg605_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg604_out,
                 Y => SharedReg605_out);

   SharedReg606_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product6_1_impl_out,
                 Y => SharedReg606_out);

   SharedReg607_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg606_out,
                 Y => SharedReg607_out);

   SharedReg608_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg607_out,
                 Y => SharedReg608_out);

   SharedReg609_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product6_2_impl_out,
                 Y => SharedReg609_out);

   SharedReg610_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg609_out,
                 Y => SharedReg610_out);

   SharedReg611_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg610_out,
                 Y => SharedReg611_out);

   SharedReg612_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product6_3_impl_out,
                 Y => SharedReg612_out);

   SharedReg613_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg612_out,
                 Y => SharedReg613_out);

   SharedReg614_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg613_out,
                 Y => SharedReg614_out);

   SharedReg615_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product6_4_impl_out,
                 Y => SharedReg615_out);

   SharedReg616_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg615_out,
                 Y => SharedReg616_out);

   SharedReg617_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg616_out,
                 Y => SharedReg617_out);

   SharedReg618_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product6_5_impl_out,
                 Y => SharedReg618_out);

   SharedReg619_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg618_out,
                 Y => SharedReg619_out);

   SharedReg620_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg619_out,
                 Y => SharedReg620_out);

   SharedReg621_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product6_6_impl_out,
                 Y => SharedReg621_out);

   SharedReg622_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg621_out,
                 Y => SharedReg622_out);

   SharedReg623_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg622_out,
                 Y => SharedReg623_out);

   SharedReg624_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product23_0_impl_out,
                 Y => SharedReg624_out);

   SharedReg625_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg624_out,
                 Y => SharedReg625_out);

   SharedReg626_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg625_out,
                 Y => SharedReg626_out);

   SharedReg627_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product23_1_impl_out,
                 Y => SharedReg627_out);

   SharedReg628_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg627_out,
                 Y => SharedReg628_out);

   SharedReg629_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg628_out,
                 Y => SharedReg629_out);

   SharedReg630_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product23_2_impl_out,
                 Y => SharedReg630_out);

   SharedReg631_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg630_out,
                 Y => SharedReg631_out);

   SharedReg632_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg631_out,
                 Y => SharedReg632_out);

   SharedReg633_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product23_3_impl_out,
                 Y => SharedReg633_out);

   SharedReg634_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg633_out,
                 Y => SharedReg634_out);

   SharedReg635_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg634_out,
                 Y => SharedReg635_out);

   SharedReg636_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product23_4_impl_out,
                 Y => SharedReg636_out);

   SharedReg637_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg636_out,
                 Y => SharedReg637_out);

   SharedReg638_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg637_out,
                 Y => SharedReg638_out);

   SharedReg639_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product23_5_impl_out,
                 Y => SharedReg639_out);

   SharedReg640_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg639_out,
                 Y => SharedReg640_out);

   SharedReg641_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg640_out,
                 Y => SharedReg641_out);

   SharedReg642_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product23_6_impl_out,
                 Y => SharedReg642_out);

   SharedReg643_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg642_out,
                 Y => SharedReg643_out);

   SharedReg644_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg643_out,
                 Y => SharedReg644_out);

   SharedReg645_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product33_0_impl_out,
                 Y => SharedReg645_out);

   SharedReg646_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg645_out,
                 Y => SharedReg646_out);

   SharedReg647_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg646_out,
                 Y => SharedReg647_out);

   SharedReg648_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product33_1_impl_out,
                 Y => SharedReg648_out);

   SharedReg649_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg648_out,
                 Y => SharedReg649_out);

   SharedReg650_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg649_out,
                 Y => SharedReg650_out);

   SharedReg651_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product33_2_impl_out,
                 Y => SharedReg651_out);

   SharedReg652_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg651_out,
                 Y => SharedReg652_out);

   SharedReg653_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg652_out,
                 Y => SharedReg653_out);

   SharedReg654_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product33_3_impl_out,
                 Y => SharedReg654_out);

   SharedReg655_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg654_out,
                 Y => SharedReg655_out);

   SharedReg656_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg655_out,
                 Y => SharedReg656_out);

   SharedReg657_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product33_4_impl_out,
                 Y => SharedReg657_out);

   SharedReg658_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg657_out,
                 Y => SharedReg658_out);

   SharedReg659_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg658_out,
                 Y => SharedReg659_out);

   SharedReg660_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product33_5_impl_out,
                 Y => SharedReg660_out);

   SharedReg661_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg660_out,
                 Y => SharedReg661_out);

   SharedReg662_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg661_out,
                 Y => SharedReg662_out);

   SharedReg663_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product33_6_impl_out,
                 Y => SharedReg663_out);

   SharedReg664_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg663_out,
                 Y => SharedReg664_out);

   SharedReg665_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg664_out,
                 Y => SharedReg665_out);

   SharedReg666_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract4_0_impl_out,
                 Y => SharedReg666_out);

   SharedReg667_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg666_out,
                 Y => SharedReg667_out);

   SharedReg668_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg667_out,
                 Y => SharedReg668_out);

   SharedReg669_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg668_out,
                 Y => SharedReg669_out);

   SharedReg670_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg669_out,
                 Y => SharedReg670_out);

   SharedReg671_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg670_out,
                 Y => SharedReg671_out);

   SharedReg672_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract4_1_impl_out,
                 Y => SharedReg672_out);

   SharedReg673_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg672_out,
                 Y => SharedReg673_out);

   SharedReg674_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg673_out,
                 Y => SharedReg674_out);

   SharedReg675_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg674_out,
                 Y => SharedReg675_out);

   SharedReg676_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg675_out,
                 Y => SharedReg676_out);

   SharedReg677_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg676_out,
                 Y => SharedReg677_out);

   SharedReg678_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract4_2_impl_out,
                 Y => SharedReg678_out);

   SharedReg679_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg678_out,
                 Y => SharedReg679_out);

   SharedReg680_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg679_out,
                 Y => SharedReg680_out);

   SharedReg681_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg680_out,
                 Y => SharedReg681_out);

   SharedReg682_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg681_out,
                 Y => SharedReg682_out);

   SharedReg683_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract4_3_impl_out,
                 Y => SharedReg683_out);

   SharedReg684_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg683_out,
                 Y => SharedReg684_out);

   SharedReg685_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg684_out,
                 Y => SharedReg685_out);

   SharedReg686_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg685_out,
                 Y => SharedReg686_out);

   SharedReg687_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg686_out,
                 Y => SharedReg687_out);

   SharedReg688_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg687_out,
                 Y => SharedReg688_out);

   SharedReg689_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract4_4_impl_out,
                 Y => SharedReg689_out);

   SharedReg690_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg689_out,
                 Y => SharedReg690_out);

   SharedReg691_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg690_out,
                 Y => SharedReg691_out);

   SharedReg692_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg691_out,
                 Y => SharedReg692_out);

   SharedReg693_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg692_out,
                 Y => SharedReg693_out);

   SharedReg694_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract4_5_impl_out,
                 Y => SharedReg694_out);

   SharedReg695_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg694_out,
                 Y => SharedReg695_out);

   SharedReg696_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg695_out,
                 Y => SharedReg696_out);

   SharedReg697_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg696_out,
                 Y => SharedReg697_out);

   SharedReg698_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg697_out,
                 Y => SharedReg698_out);

   SharedReg699_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract4_6_impl_out,
                 Y => SharedReg699_out);

   SharedReg700_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg699_out,
                 Y => SharedReg700_out);

   SharedReg701_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg700_out,
                 Y => SharedReg701_out);

   SharedReg702_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg701_out,
                 Y => SharedReg702_out);

   SharedReg703_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg702_out,
                 Y => SharedReg703_out);

   SharedReg704_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg703_out,
                 Y => SharedReg704_out);

   SharedReg705_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract5_4_impl_out,
                 Y => SharedReg705_out);

   SharedReg706_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg705_out,
                 Y => SharedReg706_out);

   SharedReg707_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg706_out,
                 Y => SharedReg707_out);

   SharedReg708_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg707_out,
                 Y => SharedReg708_out);

   SharedReg709_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg708_out,
                 Y => SharedReg709_out);

   SharedReg710_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg709_out,
                 Y => SharedReg710_out);

   SharedReg711_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg710_out,
                 Y => SharedReg711_out);

   SharedReg712_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract5_5_impl_out,
                 Y => SharedReg712_out);

   SharedReg713_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg712_out,
                 Y => SharedReg713_out);

   SharedReg714_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg713_out,
                 Y => SharedReg714_out);

   SharedReg715_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg714_out,
                 Y => SharedReg715_out);

   SharedReg716_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg715_out,
                 Y => SharedReg716_out);

   SharedReg717_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg716_out,
                 Y => SharedReg717_out);

   SharedReg718_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product26_0_impl_out,
                 Y => SharedReg718_out);

   SharedReg719_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg718_out,
                 Y => SharedReg719_out);

   SharedReg720_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg719_out,
                 Y => SharedReg720_out);

   SharedReg721_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg720_out,
                 Y => SharedReg721_out);

   SharedReg722_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product26_1_impl_out,
                 Y => SharedReg722_out);

   SharedReg723_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg722_out,
                 Y => SharedReg723_out);

   SharedReg724_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg723_out,
                 Y => SharedReg724_out);

   SharedReg725_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg724_out,
                 Y => SharedReg725_out);

   SharedReg726_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product26_2_impl_out,
                 Y => SharedReg726_out);

   SharedReg727_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg726_out,
                 Y => SharedReg727_out);

   SharedReg728_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg727_out,
                 Y => SharedReg728_out);

   SharedReg729_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg728_out,
                 Y => SharedReg729_out);

   SharedReg730_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product26_3_impl_out,
                 Y => SharedReg730_out);

   SharedReg731_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg730_out,
                 Y => SharedReg731_out);

   SharedReg732_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg731_out,
                 Y => SharedReg732_out);

   SharedReg733_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg732_out,
                 Y => SharedReg733_out);

   SharedReg734_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product26_4_impl_out,
                 Y => SharedReg734_out);

   SharedReg735_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg734_out,
                 Y => SharedReg735_out);

   SharedReg736_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg735_out,
                 Y => SharedReg736_out);

   SharedReg737_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg736_out,
                 Y => SharedReg737_out);

   SharedReg738_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product26_5_impl_out,
                 Y => SharedReg738_out);

   SharedReg739_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg738_out,
                 Y => SharedReg739_out);

   SharedReg740_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg739_out,
                 Y => SharedReg740_out);

   SharedReg741_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg740_out,
                 Y => SharedReg741_out);

   SharedReg742_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product26_6_impl_out,
                 Y => SharedReg742_out);

   SharedReg743_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg742_out,
                 Y => SharedReg743_out);

   SharedReg744_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg743_out,
                 Y => SharedReg744_out);

   SharedReg745_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg744_out,
                 Y => SharedReg745_out);

   SharedReg746_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract7_2_impl_out,
                 Y => SharedReg746_out);

   SharedReg747_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg746_out,
                 Y => SharedReg747_out);

   SharedReg748_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg747_out,
                 Y => SharedReg748_out);

   SharedReg749_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg748_out,
                 Y => SharedReg749_out);

   SharedReg750_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg749_out,
                 Y => SharedReg750_out);

   SharedReg751_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg750_out,
                 Y => SharedReg751_out);

   SharedReg752_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg751_out,
                 Y => SharedReg752_out);

   SharedReg753_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract7_3_impl_out,
                 Y => SharedReg753_out);

   SharedReg754_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg753_out,
                 Y => SharedReg754_out);

   SharedReg755_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg754_out,
                 Y => SharedReg755_out);

   SharedReg756_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg755_out,
                 Y => SharedReg756_out);

   SharedReg757_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg756_out,
                 Y => SharedReg757_out);

   SharedReg758_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract7_4_impl_out,
                 Y => SharedReg758_out);

   SharedReg759_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg758_out,
                 Y => SharedReg759_out);

   SharedReg760_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg759_out,
                 Y => SharedReg760_out);

   SharedReg761_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg760_out,
                 Y => SharedReg761_out);

   SharedReg762_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg761_out,
                 Y => SharedReg762_out);

   SharedReg763_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg762_out,
                 Y => SharedReg763_out);

   SharedReg764_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract7_5_impl_out,
                 Y => SharedReg764_out);

   SharedReg765_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg764_out,
                 Y => SharedReg765_out);

   SharedReg766_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg765_out,
                 Y => SharedReg766_out);

   SharedReg767_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg766_out,
                 Y => SharedReg767_out);

   SharedReg768_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg767_out,
                 Y => SharedReg768_out);

   SharedReg769_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg768_out,
                 Y => SharedReg769_out);

   SharedReg770_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract7_6_impl_out,
                 Y => SharedReg770_out);

   SharedReg771_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg770_out,
                 Y => SharedReg771_out);

   SharedReg772_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg771_out,
                 Y => SharedReg772_out);

   SharedReg773_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg772_out,
                 Y => SharedReg773_out);

   SharedReg774_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg773_out,
                 Y => SharedReg774_out);

   SharedReg775_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract8_1_impl_out,
                 Y => SharedReg775_out);

   SharedReg776_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg775_out,
                 Y => SharedReg776_out);

   SharedReg777_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg776_out,
                 Y => SharedReg777_out);

   SharedReg778_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg777_out,
                 Y => SharedReg778_out);

   SharedReg779_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg778_out,
                 Y => SharedReg779_out);

   SharedReg780_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg779_out,
                 Y => SharedReg780_out);

   SharedReg781_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg780_out,
                 Y => SharedReg781_out);

   SharedReg782_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg781_out,
                 Y => SharedReg782_out);

   SharedReg783_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract8_2_impl_out,
                 Y => SharedReg783_out);

   SharedReg784_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg783_out,
                 Y => SharedReg784_out);

   SharedReg785_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg784_out,
                 Y => SharedReg785_out);

   SharedReg786_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg785_out,
                 Y => SharedReg786_out);

   SharedReg787_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg786_out,
                 Y => SharedReg787_out);

   SharedReg788_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg787_out,
                 Y => SharedReg788_out);

   SharedReg789_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg788_out,
                 Y => SharedReg789_out);

   SharedReg790_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract8_4_impl_out,
                 Y => SharedReg790_out);

   SharedReg791_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg790_out,
                 Y => SharedReg791_out);

   SharedReg792_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg791_out,
                 Y => SharedReg792_out);

   SharedReg793_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg792_out,
                 Y => SharedReg793_out);

   SharedReg794_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg793_out,
                 Y => SharedReg794_out);

   SharedReg795_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract8_5_impl_out,
                 Y => SharedReg795_out);

   SharedReg796_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg795_out,
                 Y => SharedReg796_out);

   SharedReg797_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg796_out,
                 Y => SharedReg797_out);

   SharedReg798_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg797_out,
                 Y => SharedReg798_out);

   SharedReg799_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg798_out,
                 Y => SharedReg799_out);

   SharedReg800_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product18_0_impl_out,
                 Y => SharedReg800_out);

   SharedReg801_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg800_out,
                 Y => SharedReg801_out);

   SharedReg802_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg801_out,
                 Y => SharedReg802_out);

   SharedReg803_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product18_1_impl_out,
                 Y => SharedReg803_out);

   SharedReg804_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg803_out,
                 Y => SharedReg804_out);

   SharedReg805_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg804_out,
                 Y => SharedReg805_out);

   SharedReg806_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product18_2_impl_out,
                 Y => SharedReg806_out);

   SharedReg807_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg806_out,
                 Y => SharedReg807_out);

   SharedReg808_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg807_out,
                 Y => SharedReg808_out);

   SharedReg809_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product18_3_impl_out,
                 Y => SharedReg809_out);

   SharedReg810_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg809_out,
                 Y => SharedReg810_out);

   SharedReg811_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg810_out,
                 Y => SharedReg811_out);

   SharedReg812_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product18_4_impl_out,
                 Y => SharedReg812_out);

   SharedReg813_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg812_out,
                 Y => SharedReg813_out);

   SharedReg814_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg813_out,
                 Y => SharedReg814_out);

   SharedReg815_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product18_5_impl_out,
                 Y => SharedReg815_out);

   SharedReg816_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg815_out,
                 Y => SharedReg816_out);

   SharedReg817_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg816_out,
                 Y => SharedReg817_out);

   SharedReg818_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product18_6_impl_out,
                 Y => SharedReg818_out);

   SharedReg819_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg818_out,
                 Y => SharedReg819_out);

   SharedReg820_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg819_out,
                 Y => SharedReg820_out);

   SharedReg821_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product28_0_impl_out,
                 Y => SharedReg821_out);

   SharedReg822_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg821_out,
                 Y => SharedReg822_out);

   SharedReg823_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg822_out,
                 Y => SharedReg823_out);

   SharedReg824_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg823_out,
                 Y => SharedReg824_out);

   SharedReg825_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product28_1_impl_out,
                 Y => SharedReg825_out);

   SharedReg826_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg825_out,
                 Y => SharedReg826_out);

   SharedReg827_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg826_out,
                 Y => SharedReg827_out);

   SharedReg828_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg827_out,
                 Y => SharedReg828_out);

   SharedReg829_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product28_2_impl_out,
                 Y => SharedReg829_out);

   SharedReg830_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg829_out,
                 Y => SharedReg830_out);

   SharedReg831_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg830_out,
                 Y => SharedReg831_out);

   SharedReg832_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg831_out,
                 Y => SharedReg832_out);

   SharedReg833_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product28_3_impl_out,
                 Y => SharedReg833_out);

   SharedReg834_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg833_out,
                 Y => SharedReg834_out);

   SharedReg835_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg834_out,
                 Y => SharedReg835_out);

   SharedReg836_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg835_out,
                 Y => SharedReg836_out);

   SharedReg837_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product28_4_impl_out,
                 Y => SharedReg837_out);

   SharedReg838_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg837_out,
                 Y => SharedReg838_out);

   SharedReg839_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg838_out,
                 Y => SharedReg839_out);

   SharedReg840_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg839_out,
                 Y => SharedReg840_out);

   SharedReg841_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product28_5_impl_out,
                 Y => SharedReg841_out);

   SharedReg842_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg841_out,
                 Y => SharedReg842_out);

   SharedReg843_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg842_out,
                 Y => SharedReg843_out);

   SharedReg844_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg843_out,
                 Y => SharedReg844_out);

   SharedReg845_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product28_6_impl_out,
                 Y => SharedReg845_out);

   SharedReg846_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg845_out,
                 Y => SharedReg846_out);

   SharedReg847_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg846_out,
                 Y => SharedReg847_out);

   SharedReg848_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg847_out,
                 Y => SharedReg848_out);

   SharedReg849_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract9_0_impl_out,
                 Y => SharedReg849_out);

   SharedReg850_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg849_out,
                 Y => SharedReg850_out);

   SharedReg851_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg850_out,
                 Y => SharedReg851_out);

   SharedReg852_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg851_out,
                 Y => SharedReg852_out);

   SharedReg853_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg852_out,
                 Y => SharedReg853_out);

   SharedReg854_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract9_1_impl_out,
                 Y => SharedReg854_out);

   SharedReg855_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg854_out,
                 Y => SharedReg855_out);

   SharedReg856_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg855_out,
                 Y => SharedReg856_out);

   SharedReg857_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg856_out,
                 Y => SharedReg857_out);

   SharedReg858_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract9_2_impl_out,
                 Y => SharedReg858_out);

   SharedReg859_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg858_out,
                 Y => SharedReg859_out);

   SharedReg860_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg859_out,
                 Y => SharedReg860_out);

   SharedReg861_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract9_3_impl_out,
                 Y => SharedReg861_out);

   SharedReg862_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg861_out,
                 Y => SharedReg862_out);

   SharedReg863_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg862_out,
                 Y => SharedReg863_out);

   SharedReg864_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg863_out,
                 Y => SharedReg864_out);

   SharedReg865_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract9_4_impl_out,
                 Y => SharedReg865_out);

   SharedReg866_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg865_out,
                 Y => SharedReg866_out);

   SharedReg867_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg866_out,
                 Y => SharedReg867_out);

   SharedReg868_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract9_5_impl_out,
                 Y => SharedReg868_out);

   SharedReg869_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg868_out,
                 Y => SharedReg869_out);

   SharedReg870_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg869_out,
                 Y => SharedReg870_out);

   SharedReg871_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract9_6_impl_out,
                 Y => SharedReg871_out);

   SharedReg872_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg871_out,
                 Y => SharedReg872_out);

   SharedReg873_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg872_out,
                 Y => SharedReg873_out);

   SharedReg874_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg873_out,
                 Y => SharedReg874_out);

   SharedReg875_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg874_out,
                 Y => SharedReg875_out);

   SharedReg876_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract10_3_impl_out,
                 Y => SharedReg876_out);

   SharedReg877_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg876_out,
                 Y => SharedReg877_out);

   SharedReg878_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg877_out,
                 Y => SharedReg878_out);

   SharedReg879_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg878_out,
                 Y => SharedReg879_out);

   SharedReg880_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg879_out,
                 Y => SharedReg880_out);

   SharedReg881_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg880_out,
                 Y => SharedReg881_out);

   SharedReg882_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg881_out,
                 Y => SharedReg882_out);

   SharedReg883_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product50_0_impl_out,
                 Y => SharedReg883_out);

   SharedReg884_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg883_out,
                 Y => SharedReg884_out);

   SharedReg885_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg884_out,
                 Y => SharedReg885_out);

   SharedReg886_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg885_out,
                 Y => SharedReg886_out);

   SharedReg887_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product50_1_impl_out,
                 Y => SharedReg887_out);

   SharedReg888_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg887_out,
                 Y => SharedReg888_out);

   SharedReg889_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg888_out,
                 Y => SharedReg889_out);

   SharedReg890_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg889_out,
                 Y => SharedReg890_out);

   SharedReg891_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product50_2_impl_out,
                 Y => SharedReg891_out);

   SharedReg892_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg891_out,
                 Y => SharedReg892_out);

   SharedReg893_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg892_out,
                 Y => SharedReg893_out);

   SharedReg894_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg893_out,
                 Y => SharedReg894_out);

   SharedReg895_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product50_3_impl_out,
                 Y => SharedReg895_out);

   SharedReg896_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg895_out,
                 Y => SharedReg896_out);

   SharedReg897_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg896_out,
                 Y => SharedReg897_out);

   SharedReg898_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg897_out,
                 Y => SharedReg898_out);

   SharedReg899_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product50_4_impl_out,
                 Y => SharedReg899_out);

   SharedReg900_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg899_out,
                 Y => SharedReg900_out);

   SharedReg901_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg900_out,
                 Y => SharedReg901_out);

   SharedReg902_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg901_out,
                 Y => SharedReg902_out);

   SharedReg903_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product50_5_impl_out,
                 Y => SharedReg903_out);

   SharedReg904_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg903_out,
                 Y => SharedReg904_out);

   SharedReg905_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg904_out,
                 Y => SharedReg905_out);

   SharedReg906_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg905_out,
                 Y => SharedReg906_out);

   SharedReg907_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product50_6_impl_out,
                 Y => SharedReg907_out);

   SharedReg908_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg907_out,
                 Y => SharedReg908_out);

   SharedReg909_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg908_out,
                 Y => SharedReg909_out);

   SharedReg910_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg909_out,
                 Y => SharedReg910_out);

   SharedReg911_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product122_0_impl_out,
                 Y => SharedReg911_out);

   SharedReg912_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg911_out,
                 Y => SharedReg912_out);

   SharedReg913_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg912_out,
                 Y => SharedReg913_out);

   SharedReg914_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg913_out,
                 Y => SharedReg914_out);

   SharedReg915_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product122_1_impl_out,
                 Y => SharedReg915_out);

   SharedReg916_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg915_out,
                 Y => SharedReg916_out);

   SharedReg917_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg916_out,
                 Y => SharedReg917_out);

   SharedReg918_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg917_out,
                 Y => SharedReg918_out);

   SharedReg919_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product122_2_impl_out,
                 Y => SharedReg919_out);

   SharedReg920_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg919_out,
                 Y => SharedReg920_out);

   SharedReg921_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg920_out,
                 Y => SharedReg921_out);

   SharedReg922_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg921_out,
                 Y => SharedReg922_out);

   SharedReg923_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product122_3_impl_out,
                 Y => SharedReg923_out);

   SharedReg924_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg923_out,
                 Y => SharedReg924_out);

   SharedReg925_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg924_out,
                 Y => SharedReg925_out);

   SharedReg926_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg925_out,
                 Y => SharedReg926_out);

   SharedReg927_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product122_4_impl_out,
                 Y => SharedReg927_out);

   SharedReg928_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg927_out,
                 Y => SharedReg928_out);

   SharedReg929_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg928_out,
                 Y => SharedReg929_out);

   SharedReg930_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg929_out,
                 Y => SharedReg930_out);

   SharedReg931_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product122_5_impl_out,
                 Y => SharedReg931_out);

   SharedReg932_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg931_out,
                 Y => SharedReg932_out);

   SharedReg933_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg932_out,
                 Y => SharedReg933_out);

   SharedReg934_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg933_out,
                 Y => SharedReg934_out);

   SharedReg935_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product122_6_impl_out,
                 Y => SharedReg935_out);

   SharedReg936_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg935_out,
                 Y => SharedReg936_out);

   SharedReg937_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg936_out,
                 Y => SharedReg937_out);

   SharedReg938_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg937_out,
                 Y => SharedReg938_out);

   SharedReg939_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product221_0_impl_out,
                 Y => SharedReg939_out);

   SharedReg940_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg939_out,
                 Y => SharedReg940_out);

   SharedReg941_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg940_out,
                 Y => SharedReg941_out);

   SharedReg942_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product221_1_impl_out,
                 Y => SharedReg942_out);

   SharedReg943_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg942_out,
                 Y => SharedReg943_out);

   SharedReg944_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg943_out,
                 Y => SharedReg944_out);

   SharedReg945_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product221_2_impl_out,
                 Y => SharedReg945_out);

   SharedReg946_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg945_out,
                 Y => SharedReg946_out);

   SharedReg947_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg946_out,
                 Y => SharedReg947_out);

   SharedReg948_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product221_3_impl_out,
                 Y => SharedReg948_out);

   SharedReg949_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg948_out,
                 Y => SharedReg949_out);

   SharedReg950_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg949_out,
                 Y => SharedReg950_out);

   SharedReg951_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product221_4_impl_out,
                 Y => SharedReg951_out);

   SharedReg952_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg951_out,
                 Y => SharedReg952_out);

   SharedReg953_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg952_out,
                 Y => SharedReg953_out);

   SharedReg954_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product221_5_impl_out,
                 Y => SharedReg954_out);

   SharedReg955_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg954_out,
                 Y => SharedReg955_out);

   SharedReg956_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg955_out,
                 Y => SharedReg956_out);

   SharedReg957_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product221_6_impl_out,
                 Y => SharedReg957_out);

   SharedReg958_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg957_out,
                 Y => SharedReg958_out);

   SharedReg959_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg958_out,
                 Y => SharedReg959_out);

   SharedReg960_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product321_0_impl_out,
                 Y => SharedReg960_out);

   SharedReg961_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg960_out,
                 Y => SharedReg961_out);

   SharedReg962_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg961_out,
                 Y => SharedReg962_out);

   SharedReg963_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product321_1_impl_out,
                 Y => SharedReg963_out);

   SharedReg964_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg963_out,
                 Y => SharedReg964_out);

   SharedReg965_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg964_out,
                 Y => SharedReg965_out);

   SharedReg966_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product321_2_impl_out,
                 Y => SharedReg966_out);

   SharedReg967_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg966_out,
                 Y => SharedReg967_out);

   SharedReg968_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg967_out,
                 Y => SharedReg968_out);

   SharedReg969_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product321_3_impl_out,
                 Y => SharedReg969_out);

   SharedReg970_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg969_out,
                 Y => SharedReg970_out);

   SharedReg971_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg970_out,
                 Y => SharedReg971_out);

   SharedReg972_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product321_4_impl_out,
                 Y => SharedReg972_out);

   SharedReg973_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg972_out,
                 Y => SharedReg973_out);

   SharedReg974_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg973_out,
                 Y => SharedReg974_out);

   SharedReg975_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product321_5_impl_out,
                 Y => SharedReg975_out);

   SharedReg976_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg975_out,
                 Y => SharedReg976_out);

   SharedReg977_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg976_out,
                 Y => SharedReg977_out);

   SharedReg978_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product321_6_impl_out,
                 Y => SharedReg978_out);

   SharedReg979_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg978_out,
                 Y => SharedReg979_out);

   SharedReg980_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg979_out,
                 Y => SharedReg980_out);

   SharedReg981_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract23_0_impl_out,
                 Y => SharedReg981_out);

   SharedReg982_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg981_out,
                 Y => SharedReg982_out);

   SharedReg983_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg982_out,
                 Y => SharedReg983_out);

   SharedReg984_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract23_1_impl_out,
                 Y => SharedReg984_out);

   SharedReg985_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg984_out,
                 Y => SharedReg985_out);

   SharedReg986_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract23_2_impl_out,
                 Y => SharedReg986_out);

   SharedReg987_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg986_out,
                 Y => SharedReg987_out);

   SharedReg988_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg987_out,
                 Y => SharedReg988_out);

   SharedReg989_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg988_out,
                 Y => SharedReg989_out);

   SharedReg990_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract23_3_impl_out,
                 Y => SharedReg990_out);

   SharedReg991_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg990_out,
                 Y => SharedReg991_out);

   SharedReg992_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg991_out,
                 Y => SharedReg992_out);

   SharedReg993_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract23_4_impl_out,
                 Y => SharedReg993_out);

   SharedReg994_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg993_out,
                 Y => SharedReg994_out);

   SharedReg995_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg994_out,
                 Y => SharedReg995_out);

   SharedReg996_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg995_out,
                 Y => SharedReg996_out);

   SharedReg997_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract23_5_impl_out,
                 Y => SharedReg997_out);

   SharedReg998_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg997_out,
                 Y => SharedReg998_out);

   SharedReg999_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg998_out,
                 Y => SharedReg999_out);

   SharedReg1000_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg999_out,
                 Y => SharedReg1000_out);

   SharedReg1001_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract23_6_impl_out,
                 Y => SharedReg1001_out);

   SharedReg1002_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1001_out,
                 Y => SharedReg1002_out);

   SharedReg1003_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1002_out,
                 Y => SharedReg1003_out);

   SharedReg1004_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract30_0_impl_out,
                 Y => SharedReg1004_out);

   SharedReg1005_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1004_out,
                 Y => SharedReg1005_out);

   SharedReg1006_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1005_out,
                 Y => SharedReg1006_out);

   SharedReg1007_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract30_1_impl_out,
                 Y => SharedReg1007_out);

   SharedReg1008_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1007_out,
                 Y => SharedReg1008_out);

   SharedReg1009_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1008_out,
                 Y => SharedReg1009_out);

   SharedReg1010_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1009_out,
                 Y => SharedReg1010_out);

   SharedReg1011_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1010_out,
                 Y => SharedReg1011_out);

   SharedReg1012_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract30_2_impl_out,
                 Y => SharedReg1012_out);

   SharedReg1013_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1012_out,
                 Y => SharedReg1013_out);

   SharedReg1014_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1013_out,
                 Y => SharedReg1014_out);

   SharedReg1015_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1014_out,
                 Y => SharedReg1015_out);

   SharedReg1016_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1015_out,
                 Y => SharedReg1016_out);

   SharedReg1017_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract30_3_impl_out,
                 Y => SharedReg1017_out);

   SharedReg1018_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1017_out,
                 Y => SharedReg1018_out);

   SharedReg1019_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1018_out,
                 Y => SharedReg1019_out);

   SharedReg1020_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1019_out,
                 Y => SharedReg1020_out);

   SharedReg1021_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1020_out,
                 Y => SharedReg1021_out);

   SharedReg1022_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract30_4_impl_out,
                 Y => SharedReg1022_out);

   SharedReg1023_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1022_out,
                 Y => SharedReg1023_out);

   SharedReg1024_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1023_out,
                 Y => SharedReg1024_out);

   SharedReg1025_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1024_out,
                 Y => SharedReg1025_out);

   SharedReg1026_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1025_out,
                 Y => SharedReg1026_out);

   SharedReg1027_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1026_out,
                 Y => SharedReg1027_out);

   SharedReg1028_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract30_5_impl_out,
                 Y => SharedReg1028_out);

   SharedReg1029_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1028_out,
                 Y => SharedReg1029_out);

   SharedReg1030_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1029_out,
                 Y => SharedReg1030_out);

   SharedReg1031_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1030_out,
                 Y => SharedReg1031_out);

   SharedReg1032_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1031_out,
                 Y => SharedReg1032_out);

   SharedReg1033_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract30_6_impl_out,
                 Y => SharedReg1033_out);

   SharedReg1034_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1033_out,
                 Y => SharedReg1034_out);

   SharedReg1035_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1034_out,
                 Y => SharedReg1035_out);

   SharedReg1036_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1035_out,
                 Y => SharedReg1036_out);

   SharedReg1037_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract32_0_impl_out,
                 Y => SharedReg1037_out);

   SharedReg1038_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1037_out,
                 Y => SharedReg1038_out);

   SharedReg1039_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1038_out,
                 Y => SharedReg1039_out);

   SharedReg1040_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1039_out,
                 Y => SharedReg1040_out);

   SharedReg1041_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1040_out,
                 Y => SharedReg1041_out);

   SharedReg1042_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract32_1_impl_out,
                 Y => SharedReg1042_out);

   SharedReg1043_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1042_out,
                 Y => SharedReg1043_out);

   SharedReg1044_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1043_out,
                 Y => SharedReg1044_out);

   SharedReg1045_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1044_out,
                 Y => SharedReg1045_out);

   SharedReg1046_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1045_out,
                 Y => SharedReg1046_out);

   SharedReg1047_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract32_2_impl_out,
                 Y => SharedReg1047_out);

   SharedReg1048_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1047_out,
                 Y => SharedReg1048_out);

   SharedReg1049_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1048_out,
                 Y => SharedReg1049_out);

   SharedReg1050_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1049_out,
                 Y => SharedReg1050_out);

   SharedReg1051_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1050_out,
                 Y => SharedReg1051_out);

   SharedReg1052_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1051_out,
                 Y => SharedReg1052_out);

   SharedReg1053_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1052_out,
                 Y => SharedReg1053_out);

   SharedReg1054_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract32_3_impl_out,
                 Y => SharedReg1054_out);

   SharedReg1055_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1054_out,
                 Y => SharedReg1055_out);

   SharedReg1056_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1055_out,
                 Y => SharedReg1056_out);

   SharedReg1057_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1056_out,
                 Y => SharedReg1057_out);

   SharedReg1058_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1057_out,
                 Y => SharedReg1058_out);

   SharedReg1059_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1058_out,
                 Y => SharedReg1059_out);

   SharedReg1060_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract32_5_impl_out,
                 Y => SharedReg1060_out);

   SharedReg1061_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1060_out,
                 Y => SharedReg1061_out);

   SharedReg1062_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1061_out,
                 Y => SharedReg1062_out);

   SharedReg1063_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1062_out,
                 Y => SharedReg1063_out);

   SharedReg1064_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1063_out,
                 Y => SharedReg1064_out);

   SharedReg1065_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1064_out,
                 Y => SharedReg1065_out);

   SharedReg1066_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract32_6_impl_out,
                 Y => SharedReg1066_out);

   SharedReg1067_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1066_out,
                 Y => SharedReg1067_out);

   SharedReg1068_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1067_out,
                 Y => SharedReg1068_out);

   SharedReg1069_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1068_out,
                 Y => SharedReg1069_out);

   SharedReg1070_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract43_0_impl_out,
                 Y => SharedReg1070_out);

   SharedReg1071_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1070_out,
                 Y => SharedReg1071_out);

   SharedReg1072_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1071_out,
                 Y => SharedReg1072_out);

   SharedReg1073_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1072_out,
                 Y => SharedReg1073_out);

   SharedReg1074_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1073_out,
                 Y => SharedReg1074_out);

   SharedReg1075_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract44_6_impl_out,
                 Y => SharedReg1075_out);

   SharedReg1076_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1075_out,
                 Y => SharedReg1076_out);

   SharedReg1077_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1076_out,
                 Y => SharedReg1077_out);

   SharedReg1078_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1077_out,
                 Y => SharedReg1078_out);

   SharedReg1079_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1078_out,
                 Y => SharedReg1079_out);

   SharedReg1080_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1079_out,
                 Y => SharedReg1080_out);

   SharedReg1081_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract49_1_impl_out,
                 Y => SharedReg1081_out);

   SharedReg1082_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1081_out,
                 Y => SharedReg1082_out);

   SharedReg1083_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1082_out,
                 Y => SharedReg1083_out);

   SharedReg1084_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1083_out,
                 Y => SharedReg1084_out);

   SharedReg1085_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1084_out,
                 Y => SharedReg1085_out);

   SharedReg1086_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1085_out,
                 Y => SharedReg1086_out);

   SharedReg1087_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1086_out,
                 Y => SharedReg1087_out);

   SharedReg1088_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract116_6_impl_out,
                 Y => SharedReg1088_out);

   SharedReg1089_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1088_out,
                 Y => SharedReg1089_out);

   SharedReg1090_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1089_out,
                 Y => SharedReg1090_out);

   SharedReg1091_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1090_out,
                 Y => SharedReg1091_out);

   SharedReg1092_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1091_out,
                 Y => SharedReg1092_out);

   SharedReg1093_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1092_out,
                 Y => SharedReg1093_out);

   SharedReg1094_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract58_0_impl_out,
                 Y => SharedReg1094_out);

   SharedReg1095_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1094_out,
                 Y => SharedReg1095_out);

   SharedReg1096_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1095_out,
                 Y => SharedReg1096_out);

   SharedReg1097_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1096_out,
                 Y => SharedReg1097_out);

   SharedReg1098_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1097_out,
                 Y => SharedReg1098_out);

   SharedReg1099_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1098_out,
                 Y => SharedReg1099_out);

   SharedReg1100_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1099_out,
                 Y => SharedReg1100_out);

   SharedReg1101_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract125_6_impl_out,
                 Y => SharedReg1101_out);

   SharedReg1102_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1101_out,
                 Y => SharedReg1102_out);

   SharedReg1103_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant2_0_impl_out,
                 Y => SharedReg1103_out);

   SharedReg1104_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1103_out,
                 Y => SharedReg1104_out);

   SharedReg1105_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1104_out,
                 Y => SharedReg1105_out);

   SharedReg1106_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1105_out,
                 Y => SharedReg1106_out);

   SharedReg1107_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1106_out,
                 Y => SharedReg1107_out);

   SharedReg1108_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1107_out,
                 Y => SharedReg1108_out);

   SharedReg1109_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1108_out,
                 Y => SharedReg1109_out);

   SharedReg1110_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1109_out,
                 Y => SharedReg1110_out);

   SharedReg1111_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1110_out,
                 Y => SharedReg1111_out);

   SharedReg1112_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1111_out,
                 Y => SharedReg1112_out);

   SharedReg1113_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1112_out,
                 Y => SharedReg1113_out);

   SharedReg1114_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1113_out,
                 Y => SharedReg1114_out);

   SharedReg1115_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant11_0_impl_out,
                 Y => SharedReg1115_out);

   SharedReg1116_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1115_out,
                 Y => SharedReg1116_out);

   SharedReg1117_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1116_out,
                 Y => SharedReg1117_out);

   SharedReg1118_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1117_out,
                 Y => SharedReg1118_out);

   SharedReg1119_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1118_out,
                 Y => SharedReg1119_out);

   SharedReg1120_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1119_out,
                 Y => SharedReg1120_out);

   SharedReg1121_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1120_out,
                 Y => SharedReg1121_out);

   SharedReg1122_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1121_out,
                 Y => SharedReg1122_out);

   SharedReg1123_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1122_out,
                 Y => SharedReg1123_out);

   SharedReg1124_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1123_out,
                 Y => SharedReg1124_out);

   SharedReg1125_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1124_out,
                 Y => SharedReg1125_out);

   SharedReg1126_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1125_out,
                 Y => SharedReg1126_out);

   SharedReg1127_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant4_0_impl_out,
                 Y => SharedReg1127_out);

   SharedReg1128_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1127_out,
                 Y => SharedReg1128_out);

   SharedReg1129_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1128_out,
                 Y => SharedReg1129_out);

   SharedReg1130_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant13_0_impl_out,
                 Y => SharedReg1130_out);

   SharedReg1131_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1130_out,
                 Y => SharedReg1131_out);

   SharedReg1132_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant5_0_impl_out,
                 Y => SharedReg1132_out);

   SharedReg1133_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant14_0_impl_out,
                 Y => SharedReg1133_out);

   SharedReg1134_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant6_0_impl_out,
                 Y => SharedReg1134_out);

   SharedReg1135_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1134_out,
                 Y => SharedReg1135_out);

   SharedReg1136_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1135_out,
                 Y => SharedReg1136_out);

   SharedReg1137_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1136_out,
                 Y => SharedReg1137_out);

   SharedReg1138_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant15_0_impl_out,
                 Y => SharedReg1138_out);

   SharedReg1139_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1138_out,
                 Y => SharedReg1139_out);

   SharedReg1140_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1139_out,
                 Y => SharedReg1140_out);

   SharedReg1141_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1140_out,
                 Y => SharedReg1141_out);

   SharedReg1142_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant7_0_impl_out,
                 Y => SharedReg1142_out);

   SharedReg1143_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1142_out,
                 Y => SharedReg1143_out);

   SharedReg1144_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant16_0_impl_out,
                 Y => SharedReg1144_out);

   SharedReg1145_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1144_out,
                 Y => SharedReg1145_out);

   SharedReg1146_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant8_0_impl_out,
                 Y => SharedReg1146_out);

   SharedReg1147_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1146_out,
                 Y => SharedReg1147_out);

   SharedReg1148_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1147_out,
                 Y => SharedReg1148_out);

   SharedReg1149_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1148_out,
                 Y => SharedReg1149_out);

   SharedReg1150_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant17_0_impl_out,
                 Y => SharedReg1150_out);

   SharedReg1151_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1150_out,
                 Y => SharedReg1151_out);

   SharedReg1152_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1151_out,
                 Y => SharedReg1152_out);

   SharedReg1153_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1152_out,
                 Y => SharedReg1153_out);

   SharedReg1154_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant9_0_impl_out,
                 Y => SharedReg1154_out);

   SharedReg1155_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1154_out,
                 Y => SharedReg1155_out);

   SharedReg1156_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant18_0_impl_out,
                 Y => SharedReg1156_out);

   SharedReg1157_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1156_out,
                 Y => SharedReg1157_out);

   SharedReg1158_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant_0_impl_out,
                 Y => SharedReg1158_out);

   SharedReg1159_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant1_0_impl_out,
                 Y => SharedReg1159_out);
end architecture;

